`timescale 1 ns/100 ps
// Version: v11.6 SP1 11.6.1.6


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module dds(
       dds_sin,
       dds_cos,
       dac_count,
       BW_clk_c
    );
output [7:0] dds_sin;
output [7:0] dds_cos;
input  [7:1] dac_count;
input  BW_clk_c;

    wire VCC_net_1, N_130_i, GND_net_1, m131, N_134_i, N_136_i, 
        N_138_i, N_140_i, N_142_i, N_144_i, m17, m45, m71_ns, m90, 
        m105, m118, N_126_i, m128, m106, m69, m50, m133_ns_1, 
        m97_1_2_1, m97_1_2, m94, m91, m97, m73, m76, m76_1_1, m76_0, 
        m19, m74, m21, m24_1_2, m24, m14, m22, m66, m67, m69_1_2, m64, 
        m50_1, m50_1_0, m28, m2, m63_ns_1, m63_ns, m78, m84_ns_1, 
        i3_mux_7, m16_ns_1, m16_ns, i3_mux_8, m57_ns, m71_ns_1, m44_bm, 
        m44_am, m44_ns, m130_bm, m130_am, m130_ns, m136_bm, m136_am, 
        m136_ns, m9_bm, m9_am, m9_ns, m31_bm, m31_am, m31_ns, m53, 
        i2_mux_1, m86, m87, m88_ns, m100, m103, m104_ns, i3_mux_6, 
        m81_ns, m112, m109, m48, m46, m29, N_146_mux, i4_mux_0, i4_mux, 
        m102, m98, m37, m35, m140, m124, N_147_mux, m115, i5_mux, m116, 
        i4_mux_5, m138, m134, m117, m89, m32;
    
    SLE \sin_o_2_0_dreg[0]  (.D(m17), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[0]));
    CFG3 #( .INIT(8'hB8) )  \sin_o_2_0_15_0_.m138  (.A(m115), .B(
        dac_count[7]), .C(m116), .Y(m138));
    CFG3 #( .INIT(8'hD8) )  \sin_o_2_0_15_0_.m130_ns  (.A(dac_count[7])
        , .B(m130_bm), .C(m130_am), .Y(m130_ns));
    SLE \sin_o_2_0_dreg[9]  (.D(m131), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_sin[1]));
    CFG3 #( .INIT(8'h46) )  \sin_o_2_0_15_0_.m128  (.A(dac_count[6]), 
        .B(dac_count[7]), .C(N_146_mux), .Y(m128));
    SLE \sin_o_2_0_dreg[7]  (.D(m128), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[7]));
    SLE \sin_o_2_0_dreg[1]  (.D(m45), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[1]));
    CFG4 #( .INIT(16'h2760) )  \sin_o_2_0_15_0_.m63_ns_1  (.A(
        dac_count[2]), .B(dac_count[4]), .C(dac_count[5]), .D(
        dac_count[3]), .Y(m63_ns_1));
    CFG3 #( .INIT(8'h8C) )  \sin_o_2_0_15_0_.N_144_i  (.A(dac_count[6])
        , .B(dac_count[7]), .C(N_146_mux), .Y(N_144_i));
    CFG3 #( .INIT(8'h6B) )  \sin_o_2_0_15_0_.m64  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m64));
    CFG3 #( .INIT(8'h07) )  \sin_o_2_0_15_0_.m46  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m46));
    CFG3 #( .INIT(8'hB1) )  \sin_o_2_0_15_0_.m17  (.A(dac_count[6]), 
        .B(m9_ns), .C(m16_ns), .Y(m17));
    CFG3 #( .INIT(8'h38) )  \sin_o_2_0_15_0_.m19  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m19));
    CFG4 #( .INIT(16'h0C6C) )  \sin_o_2_0_15_0_.m37  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(m37));
    CFG4 #( .INIT(16'h4051) )  \sin_o_2_0_15_0_.m115  (.A(dac_count[5])
        , .B(dac_count[4]), .C(m46), .D(m112), .Y(m115));
    CFG4 #( .INIT(16'hC318) )  \sin_o_2_0_15_0_.m86  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(m86));
    CFG3 #( .INIT(8'h7C) )  \sin_o_2_0_15_0_.m78  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m78));
    CFG4 #( .INIT(16'hB60E) )  \sin_o_2_0_15_0_.m63_ns  (.A(
        dac_count[1]), .B(dac_count[3]), .C(dac_count[5]), .D(m63_ns_1)
        , .Y(m63_ns));
    CFG3 #( .INIT(8'h62) )  \sin_o_2_0_15_0_.m29  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m29));
    CFG4 #( .INIT(16'h3323) )  \sin_o_2_0_15_0_.m120  (.A(dac_count[4])
        , .B(dac_count[7]), .C(m46), .D(dac_count[5]), .Y(N_147_mux));
    SLE \sin_o_2_0_dreg[6]  (.D(N_126_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_cos[6]));
    CFG3 #( .INIT(8'h1D) )  \sin_o_2_0_15_0_.m108  (.A(m106), .B(
        dac_count[7]), .C(m109), .Y(i5_mux));
    CFG4 #( .INIT(16'h5D19) )  \sin_o_2_0_15_0_.m133_ns_1  (.A(
        dac_count[6]), .B(dac_count[7]), .C(m57_ns), .D(m63_ns), .Y(
        m133_ns_1));
    SLE \sin_o_2_0_dreg[8]  (.D(N_130_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[0]));
    CFG3 #( .INIT(8'h72) )  \sin_o_2_0_15_0_.N_130_i  (.A(dac_count[6])
        , .B(m9_ns), .C(m16_ns), .Y(N_130_i));
    VCC VCC (.Y(VCC_net_1));
    SLE \sin_o_2_0_dreg[11]  (.D(N_136_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[3]));
    CFG4 #( .INIT(16'h1F10) )  \sin_o_2_0_15_0_.m98  (.A(dac_count[2]), 
        .B(dac_count[3]), .C(dac_count[5]), .D(m67), .Y(m98));
    CFG4 #( .INIT(16'h7F70) )  \sin_o_2_0_15_0_.m91  (.A(dac_count[2]), 
        .B(dac_count[3]), .C(dac_count[5]), .D(m46), .Y(m91));
    CFG4 #( .INIT(16'hD1F3) )  \sin_o_2_0_15_0_.m140  (.A(dac_count[4])
        , .B(dac_count[7]), .C(N_146_mux), .D(m109), .Y(m140));
    CFG3 #( .INIT(8'h78) )  \sin_o_2_0_15_0_.m73  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m73));
    CFG3 #( .INIT(8'h8B) )  \sin_o_2_0_15_0_.m136_am  (.A(m91), .B(
        dac_count[4]), .C(m102), .Y(m136_am));
    CFG3 #( .INIT(8'h39) )  \sin_o_2_0_15_0_.m84_ns_1  (.A(
        dac_count[1]), .B(dac_count[2]), .C(dac_count[3]), .Y(m84_ns_1)
        );
    SLE \sin_o_2_0_dreg[4]  (.D(m105), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[4]));
    CFG3 #( .INIT(8'h47) )  \sin_o_2_0_15_0_.N_126_i  (.A(m124), .B(
        dac_count[6]), .C(N_147_mux), .Y(N_126_i));
    CFG3 #( .INIT(8'hC7) )  \sin_o_2_0_15_0_.m87  (.A(dac_count[3]), 
        .B(dac_count[5]), .C(m19), .Y(m87));
    CFG4 #( .INIT(16'hD782) )  \sin_o_2_0_15_0_.m16_ns  (.A(
        dac_count[4]), .B(dac_count[5]), .C(m14), .D(m16_ns_1), .Y(
        m16_ns));
    CFG4 #( .INIT(16'h5702) )  \sin_o_2_0_15_0_.m100  (.A(dac_count[4])
        , .B(dac_count[5]), .C(m46), .D(m98), .Y(m100));
    CFG3 #( .INIT(8'hB8) )  \sin_o_2_0_15_0_.m89  (.A(m88_ns), .B(
        dac_count[7]), .C(i3_mux_7), .Y(m89));
    CFG3 #( .INIT(8'hD1) )  \sin_o_2_0_15_0_.m44_am  (.A(m35), .B(
        dac_count[4]), .C(m37), .Y(m44_am));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m134  (.A(m88_ns), .B(
        dac_count[7]), .C(i3_mux_7), .Y(m134));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m130_am  (.A(i4_mux), .B(
        dac_count[5]), .C(i4_mux_0), .Y(m130_am));
    CFG3 #( .INIT(8'h31) )  \sin_o_2_0_15_0_.m74  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m74));
    CFG3 #( .INIT(8'h34) )  \sin_o_2_0_15_0_.m66  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m66));
    CFG4 #( .INIT(16'h74FC) )  \sin_o_2_0_15_0_.m124  (.A(dac_count[4])
        , .B(dac_count[7]), .C(N_146_mux), .D(m109), .Y(m124));
    CFG4 #( .INIT(16'h3D0F) )  \sin_o_2_0_15_0_.m97_1_2  (.A(
        dac_count[3]), .B(m97_1_2_1), .C(dac_count[7]), .D(
        dac_count[4]), .Y(m97_1_2));
    CFG3 #( .INIT(8'hD1) )  \sin_o_2_0_15_0_.m130_bm  (.A(m35), .B(
        dac_count[4]), .C(m37), .Y(m130_bm));
    CFG3 #( .INIT(8'h74) )  \sin_o_2_0_15_0_.N_136_i  (.A(m81_ns), .B(
        dac_count[6]), .C(m134), .Y(N_136_i));
    CFG4 #( .INIT(16'h497F) )  \sin_o_2_0_15_0_.m53  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(m53));
    CFG3 #( .INIT(8'hB1) )  \sin_o_2_0_15_0_.m105  (.A(dac_count[6]), 
        .B(m97), .C(m104_ns), .Y(m105));
    CFG3 #( .INIT(8'h72) )  \sin_o_2_0_15_0_.N_138_i  (.A(dac_count[6])
        , .B(m97), .C(m136_ns), .Y(N_138_i));
    CFG3 #( .INIT(8'h70) )  \sin_o_2_0_15_0_.m94  (.A(dac_count[2]), 
        .B(dac_count[3]), .C(dac_count[5]), .Y(m94));
    CFG3 #( .INIT(8'hE4) )  \sin_o_2_0_15_0_.m116  (.A(dac_count[4]), 
        .B(dac_count[5]), .C(m106), .Y(m116));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h01) )  \sin_o_2_0_15_0_.m50_0  (.A(dac_count[4]), 
        .B(dac_count[5]), .C(m46), .Y(m76));
    SLE \sin_o_2_0_dreg[13]  (.D(N_140_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[5]));
    CFG3 #( .INIT(8'hB8) )  \sin_o_2_0_15_0_.m44_ns  (.A(m44_bm), .B(
        dac_count[7]), .C(m44_am), .Y(m44_ns));
    CFG3 #( .INIT(8'hD1) )  \sin_o_2_0_15_0_.m90  (.A(m81_ns), .B(
        dac_count[6]), .C(m89), .Y(m90));
    CFG4 #( .INIT(16'h11CF) )  \sin_o_2_0_15_0_.m69_1_2  (.A(
        dac_count[2]), .B(dac_count[4]), .C(m64), .D(dac_count[5]), .Y(
        m69_1_2));
    CFG4 #( .INIT(16'h139B) )  \sin_o_2_0_15_0_.m71_ns_1  (.A(
        dac_count[6]), .B(dac_count[7]), .C(m63_ns), .D(m69), .Y(
        m71_ns_1));
    CFG3 #( .INIT(8'h3E) )  \sin_o_2_0_15_0_.m67  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m67));
    CFG4 #( .INIT(16'hEE50) )  \sin_o_2_0_15_0_.N_134_i  (.A(
        dac_count[7]), .B(m69), .C(m50), .D(m133_ns_1), .Y(N_134_i));
    CFG4 #( .INIT(16'hDDA0) )  \sin_o_2_0_15_0_.m69  (.A(dac_count[4]), 
        .B(m66), .C(m67), .D(m69_1_2), .Y(m69));
    CFG3 #( .INIT(8'h52) )  \sin_o_2_0_15_0_.m28  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m28));
    CFG4 #( .INIT(16'hFFCE) )  \sin_o_2_0_15_0_.m50  (.A(dac_count[5]), 
        .B(m50_1), .C(m50_1_0), .D(m76), .Y(m50));
    CFG3 #( .INIT(8'h54) )  \sin_o_2_0_15_0_.m21  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m21));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m117  (.A(m115), .B(
        dac_count[7]), .C(m116), .Y(m117));
    CFG3 #( .INIT(8'h80) )  \sin_o_2_0_15_0_.m109  (.A(dac_count[2]), 
        .B(dac_count[3]), .C(dac_count[5]), .Y(m109));
    CFG4 #( .INIT(16'h0F02) )  \sin_o_2_0_15_0_.m76  (.A(m73), .B(
        dac_count[5]), .C(m76), .D(m76_1_1), .Y(m76_0));
    CFG4 #( .INIT(16'h72D8) )  \sin_o_2_0_15_0_.m111  (.A(dac_count[4])
        , .B(dac_count[7]), .C(i5_mux), .D(dac_count[5]), .Y(i4_mux_5));
    CFG4 #( .INIT(16'h6A73) )  \sin_o_2_0_15_0_.m35  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(m35));
    CFG3 #( .INIT(8'hB8) )  \sin_o_2_0_15_0_.m136_ns  (.A(m136_bm), .B(
        dac_count[7]), .C(m136_am), .Y(m136_ns));
    CFG3 #( .INIT(8'hD1) )  \sin_o_2_0_15_0_.m32  (.A(m24), .B(
        dac_count[7]), .C(m31_ns), .Y(m32));
    CFG3 #( .INIT(8'h39) )  \sin_o_2_0_15_0_.m22  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m22));
    CFG4 #( .INIT(16'h3FF8) )  \sin_o_2_0_15_0_.m106  (.A(dac_count[1])
        , .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(
        m106));
    SLE \sin_o_2_0_dreg[3]  (.D(m90), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[3]));
    CFG3 #( .INIT(8'h67) )  \sin_o_2_0_15_0_.m48  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m48));
    SLE \sin_o_2_0_dreg[5]  (.D(m118), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[5]));
    SLE \sin_o_2_0_dreg[2]  (.D(m71_ns), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dds_cos[2]));
    CFG3 #( .INIT(8'h35) )  \sin_o_2_0_15_0_.m14  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m14));
    CFG3 #( .INIT(8'hB8) )  \sin_o_2_0_15_0_.m131  (.A(m32), .B(
        dac_count[6]), .C(m130_ns), .Y(m131));
    CFG3 #( .INIT(8'h01) )  \sin_o_2_0_15_0_.m112  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .Y(m112));
    CFG4 #( .INIT(16'h6431) )  \sin_o_2_0_15_0_.m84_ns  (.A(
        dac_count[5]), .B(dac_count[4]), .C(m78), .D(m84_ns_1), .Y(
        i3_mux_7));
    CFG3 #( .INIT(8'hB8) )  \sin_o_2_0_15_0_.m31_ns  (.A(m31_bm), .B(
        dac_count[4]), .C(m31_am), .Y(m31_ns));
    CFG4 #( .INIT(16'h02F7) )  \sin_o_2_0_15_0_.m16_ns_1  (.A(
        dac_count[1]), .B(dac_count[3]), .C(dac_count[5]), .D(i3_mux_8)
        , .Y(m16_ns_1));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m81_ns  (.A(m76_0), .B(
        dac_count[7]), .C(i3_mux_6), .Y(m81_ns));
    CFG4 #( .INIT(16'h4B9C) )  \sin_o_2_0_15_0_.m56  (.A(dac_count[1]), 
        .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(
        i2_mux_1));
    CFG4 #( .INIT(16'h05EE) )  \sin_o_2_0_15_0_.m24  (.A(dac_count[5]), 
        .B(m21), .C(m19), .D(m24_1_2), .Y(m24));
    CFG3 #( .INIT(8'hE4) )  \sin_o_2_0_15_0_.m88_ns  (.A(dac_count[4]), 
        .B(m86), .C(m87), .Y(m88_ns));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m45  (.A(m32), .B(
        dac_count[6]), .C(m44_ns), .Y(m45));
    CFG3 #( .INIT(8'h1D) )  \sin_o_2_0_15_0_.N_142_i  (.A(m140), .B(
        dac_count[6]), .C(N_147_mux), .Y(N_142_i));
    CFG3 #( .INIT(8'h2E) )  \sin_o_2_0_15_0_.N_140_i  (.A(m138), .B(
        dac_count[6]), .C(i4_mux_5), .Y(N_140_i));
    CFG4 #( .INIT(16'h5B06) )  \sin_o_2_0_15_0_.m9_bm  (.A(
        dac_count[1]), .B(dac_count[2]), .C(dac_count[3]), .D(
        dac_count[5]), .Y(m9_bm));
    CFG4 #( .INIT(16'h5702) )  \sin_o_2_0_15_0_.m136_bm  (.A(
        dac_count[4]), .B(dac_count[5]), .C(m46), .D(m98), .Y(m136_bm));
    CFG3 #( .INIT(8'hCA) )  \sin_o_2_0_15_0_.m42  (.A(dac_count[1]), 
        .B(m22), .C(dac_count[4]), .Y(i4_mux_0));
    CFG3 #( .INIT(8'h10) )  \sin_o_2_0_15_0_.m122  (.A(dac_count[4]), 
        .B(dac_count[5]), .C(m112), .Y(N_146_mux));
    CFG3 #( .INIT(8'h87) )  \sin_o_2_0_15_0_.m12x  (.A(dac_count[2]), 
        .B(dac_count[3]), .C(dac_count[5]), .Y(i3_mux_8));
    CFG3 #( .INIT(8'hE4) )  \sin_o_2_0_15_0_.m57_ns  (.A(dac_count[4]), 
        .B(m53), .C(i2_mux_1), .Y(m57_ns));
    CFG3 #( .INIT(8'h02) )  \sin_o_2_0_15_0_.m50_2  (.A(dac_count[4]), 
        .B(dac_count[5]), .C(m48), .Y(m50_1));
    CFG4 #( .INIT(16'h30DD) )  \sin_o_2_0_15_0_.m97  (.A(m94), .B(
        dac_count[4]), .C(m91), .D(m97_1_2), .Y(m97));
    SLE \sin_o_2_0_dreg[15]  (.D(N_144_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[7]));
    SLE \sin_o_2_0_dreg[14]  (.D(N_142_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[6]));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m44_bm  (.A(i4_mux), .B(
        dac_count[5]), .C(i4_mux_0), .Y(m44_bm));
    CFG2 #( .INIT(4'h4) )  \sin_o_2_0_15_0_.m2  (.A(dac_count[3]), .B(
        dac_count[2]), .Y(m2));
    CFG3 #( .INIT(8'h8B) )  \sin_o_2_0_15_0_.m103  (.A(m91), .B(
        dac_count[4]), .C(m102), .Y(m103));
    CFG4 #( .INIT(16'h58A7) )  \sin_o_2_0_15_0_.m9_am  (.A(
        dac_count[1]), .B(dac_count[2]), .C(dac_count[3]), .D(
        dac_count[5]), .Y(m9_am));
    CFG4 #( .INIT(16'h31B9) )  \sin_o_2_0_15_0_.m76_1_1  (.A(
        dac_count[5]), .B(dac_count[4]), .C(m19), .D(m74), .Y(m76_1_1));
    CFG3 #( .INIT(8'hD8) )  \sin_o_2_0_15_0_.m9_ns  (.A(dac_count[4]), 
        .B(m9_bm), .C(m9_am), .Y(m9_ns));
    CFG4 #( .INIT(16'h159D) )  \sin_o_2_0_15_0_.m24_1_2  (.A(
        dac_count[4]), .B(dac_count[5]), .C(m14), .D(m22), .Y(m24_1_2));
    SLE \sin_o_2_0_dreg[12]  (.D(N_138_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[4]));
    CFG4 #( .INIT(16'h478B) )  \sin_o_2_0_15_0_.m40  (.A(dac_count[1]), 
        .B(dac_count[4]), .C(m22), .D(m2), .Y(i4_mux));
    CFG3 #( .INIT(8'h8B) )  \sin_o_2_0_15_0_.m118  (.A(m117), .B(
        dac_count[6]), .C(i4_mux_5), .Y(m118));
    CFG4 #( .INIT(16'h031F) )  \sin_o_2_0_15_0_.m102  (.A(dac_count[1])
        , .B(dac_count[2]), .C(dac_count[3]), .D(dac_count[5]), .Y(
        m102));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m31_bm  (.A(m28), .B(
        dac_count[5]), .C(m29), .Y(m31_bm));
    CFG4 #( .INIT(16'h077F) )  \sin_o_2_0_15_0_.m97_1_2_1  (.A(
        dac_count[1]), .B(dac_count[2]), .C(dac_count[3]), .D(
        dac_count[5]), .Y(m97_1_2_1));
    CFG4 #( .INIT(16'h1D2E) )  \sin_o_2_0_15_0_.m50_1_0  (.A(
        dac_count[1]), .B(dac_count[4]), .C(m28), .D(m2), .Y(m50_1_0));
    CFG3 #( .INIT(8'hE2) )  \sin_o_2_0_15_0_.m104_ns  (.A(m100), .B(
        dac_count[7]), .C(m103), .Y(m104_ns));
    SLE \sin_o_2_0_dreg[10]  (.D(N_134_i), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dds_sin[2]));
    CFG4 #( .INIT(16'h50BB) )  \sin_o_2_0_15_0_.m71_ns  (.A(
        dac_count[6]), .B(m57_ns), .C(m50), .D(m71_ns_1), .Y(m71_ns));
    CFG4 #( .INIT(16'h93D7) )  \sin_o_2_0_15_0_.m80  (.A(dac_count[5]), 
        .B(dac_count[4]), .C(m19), .D(m78), .Y(i3_mux_6));
    CFG4 #( .INIT(16'h6D60) )  \sin_o_2_0_15_0_.m31_am  (.A(
        dac_count[1]), .B(dac_count[2]), .C(dac_count[3]), .D(
        dac_count[5]), .Y(m31_am));
    
endmodule


module led_igloo(
       sdv_count,
       temp_count_data,
       BW_c,
       fpga_shift_2,
       BW_out_c,
       fpga_count,
       \data_from_adc[6] ,
       \data_from_adc[7] ,
       \data_from_adc[8] ,
       fr_adc_count,
       temp3,
       dac1_db_c,
       \data_from_adc[0] ,
       \data_from_adc[1] ,
       \data_from_adc[3] ,
       \data_from_adc[2] ,
       \data_from_adc[4] ,
       \data_from_adc[5] ,
       temp1,
       temp2,
       SENSE_DOUT_c,
       dac_count,
       temp_count,
       dds_cos,
       dds_sin,
       adc_d0_c,
       freq_10,
       freq_11,
       freq_0,
       freq_1,
       freq_13,
       freq_14,
       freq_15,
       freq_6,
       freq_2,
       temp_sck_c,
       BW_clk_c_i_0,
       BW_clk_c,
       GPIO4_c,
       temp_sck_c_i_0,
       temp_so_c,
       dac1_clk_c,
       SENSE_CS_1_c,
       GPIO16_c,
       clk_dac2,
       GPIO14_c,
       GPIO7_c,
       temp3_csn_c,
       temp2_csn_c,
       temp1_csn_c,
       GPIO11_c,
       oclk_1_c,
       GPIO10_c,
       dac2_clk_c,
       adc_of_c,
       adc_oen_c,
       adc_clk_c,
       GPS_I1_c,
       GPS_I0_c,
       GPS2_Q1_c,
       GPS2_Q0_c,
       GPS2_LD_c,
       GPS1_Q1_c,
       GPS1_Q0_c,
       GPS1_LD_c,
       GPS1_I1_c,
       GPS1_I0_c,
       GPIO9_c,
       GPIO6_c,
       osc_vcc_c,
       ANTF_n2_c,
       ANTF_n1_c,
       GPIO3_c,
       GPIO5_c
    );
output [1:0] sdv_count;
output [4:0] temp_count_data;
input  [14:0] BW_c;
output [14:0] fpga_shift_2;
output [14:0] BW_out_c;
output [14:0] fpga_count;
output [11:0] \data_from_adc[6] ;
output [11:0] \data_from_adc[7] ;
output [11:0] \data_from_adc[8] ;
output [3:1] fr_adc_count;
output [15:0] temp3;
output [13:5] dac1_db_c;
output [11:0] \data_from_adc[0] ;
output [11:0] \data_from_adc[1] ;
output [11:0] \data_from_adc[3] ;
output [11:0] \data_from_adc[2] ;
output [11:0] \data_from_adc[4] ;
output [11:0] \data_from_adc[5] ;
output [15:0] temp1;
output [15:0] temp2;
output [1:1] SENSE_DOUT_c;
output [7:1] dac_count;
output [31:0] temp_count;
output [7:0] dds_cos;
output [7:0] dds_sin;
input  [13:0] adc_d0_c;
output freq_10;
output freq_11;
output freq_0;
output freq_1;
output freq_13;
output freq_14;
output freq_15;
output freq_6;
output freq_2;
input  temp_sck_c;
input  BW_clk_c_i_0;
input  BW_clk_c;
input  GPIO4_c;
input  temp_sck_c_i_0;
input  temp_so_c;
output dac1_clk_c;
output SENSE_CS_1_c;
output GPIO16_c;
output clk_dac2;
output GPIO14_c;
output GPIO7_c;
output temp3_csn_c;
output temp2_csn_c;
output temp1_csn_c;
input  GPIO11_c;
output oclk_1_c;
input  GPIO10_c;
output dac2_clk_c;
input  adc_of_c;
input  adc_oen_c;
input  adc_clk_c;
input  GPS_I1_c;
input  GPS_I0_c;
input  GPS2_Q1_c;
input  GPS2_Q0_c;
input  GPS2_LD_c;
input  GPS1_Q1_c;
input  GPS1_Q0_c;
input  GPS1_LD_c;
input  GPS1_I1_c;
input  GPS1_I0_c;
input  GPIO9_c;
input  GPIO6_c;
input  osc_vcc_c;
input  ANTF_n2_c;
input  ANTF_n1_c;
output GPIO3_c;
output GPIO5_c;

    wire \fpga_count_s[0] , \cnt_freq[0]_net_1 , \cnt_freq_s[0] , 
        \temp_state[1]_net_1 , \temp_state_i_0[1] , 
        \temp_state[0]_net_1 , \temp_state_i_0[0] , \sdv_count_i_0[1] , 
        \sdv_count_i_0[0] , temp_state26, N_449_i, fpga_flag_net_1, 
        fpga_flag_i, VCC_net_1, N_9_i_0, un1_temp_state28_0_net_1, 
        GND_net_1, N_7_i_0, N_28_i_0, N_11_i_0, N_33, 
        \fpga_data_receive[3]_net_1 , \fpga_data_receive[4]_net_1 , 
        \fpga_data_receive[5]_net_1 , \fpga_data_receive[6]_net_1 , 
        \fpga_data_receive[7]_net_1 , \fpga_data_receive[8]_net_1 , 
        \fpga_data_receive[9]_net_1 , \fpga_data_receive[10]_net_1 , 
        \fpga_data_receive[11]_net_1 , \fpga_data_receive[12]_net_1 , 
        \fpga_data_receive[13]_net_1 , \fpga_data_receive[14]_net_1 , 
        \fpga_data_receive[0]_net_1 , \fpga_data_receive[1]_net_1 , 
        \fpga_data_receive[2]_net_1 , N_11_i_0_0, 
        \temp_state[2]_net_1 , \temp_state_7[2] , \sdv_count_1[1] , 
        \temp_state_7[0] , \data_from_adc[7]_163 , 
        \data_from_adc[7]_164 , \data_from_adc[6]_141 , 
        \data_from_adc[6]_142 , \data_from_adc[6]_143 , 
        \data_from_adc[6]_144 , \data_from_adc[6]_145 , 
        \data_from_adc[6]_146 , \data_from_adc[6]_147 , 
        \data_from_adc[6]_148 , \data_from_adc[6]_149 , 
        \data_from_adc[6]_150 , \data_from_adc[6]_151 , 
        \data_from_adc[6]_152 , \data_from_adc[8]_172 , 
        \data_from_adc[8]_173 , \data_from_adc[8]_174 , 
        \data_from_adc[8]_175 , \data_from_adc[8]_176 , 
        \data_from_adc[7]_153 , \data_from_adc[7]_154 , 
        \data_from_adc[7]_155 , \data_from_adc[7]_156 , 
        \data_from_adc[7]_157 , \data_from_adc[7]_158 , 
        \data_from_adc[7]_159 , \data_from_adc[7]_160 , 
        \data_from_adc[7]_161 , \data_from_adc[7]_162 , 
        \state[1]_net_1 , N_40_i_0, un1_state15_0_net_1, freq3_i_0, 
        \un1_data_from_adc[2]_1_i_i_0 , \un1_data_from_adc[2]_2 , 
        freq9_net_1, freq3, \data_from_adc[8]_165 , 
        \data_from_adc[8]_166 , \data_from_adc[8]_167 , 
        \data_from_adc[8]_168 , \data_from_adc[8]_169 , 
        \data_from_adc[8]_170 , \data_from_adc[8]_171 , temp3_43, 
        temp3_44, temp3_45, temp3_46, temp3_47, temp3_48, temp3_49, 
        freq15_i_0, \fr_adc_count_5_i_0[2] , 
        \un1_data_from_adc[2]_i_0 , \fr_adc_count_5[1] , 
        \fr_adc_count_5[2] , freq9_i_0_net_1, \state[0]_net_1 , N_42, 
        temp3_34, temp3_35, temp3_36, temp3_37, temp3_38, temp3_39, 
        temp3_40, temp3_41, temp3_42, \data_from_adc[0]_77 , 
        \data_from_adc[0]_78 , \data_from_adc[0]_79 , 
        \data_from_adc[0]_80 , dac1_db_8_306_i_m2_net_1, 
        dac1_db_8_0_296_i_m2_net_1, dac1_db_8_1_286_i_m2_net_1, 
        dac1_db_8_2_276_i_m2_net_1, dac1_db_8_3_266_i_m2_net_1, 
        dac1_db_8_4_256_i_m2_net_1, dac1_db_8_5_246_i_m2_net_1, 
        dac1_db_8_6_236_i_m2_net_1, dac1_db_0_sqmuxa_net_1, 
        \data_from_adc[1]_86 , \data_from_adc[1]_87 , 
        \data_from_adc[1]_88 , \data_from_adc[1]_89 , 
        \data_from_adc[1]_90 , \data_from_adc[1]_91 , 
        \data_from_adc[1]_92 , \data_from_adc[0]_69 , 
        \data_from_adc[0]_70 , \data_from_adc[0]_71 , 
        \data_from_adc[0]_72 , \data_from_adc[0]_73 , 
        \data_from_adc[0]_74 , \data_from_adc[0]_75 , 
        \data_from_adc[0]_76 , \data_from_adc[2]_95 , 
        \data_from_adc[2]_96 , \data_from_adc[2]_97 , 
        \data_from_adc[2]_98 , \data_from_adc[2]_99 , 
        \data_from_adc[2]_100 , \data_from_adc[2]_101 , 
        \data_from_adc[2]_102 , \data_from_adc[2]_103 , 
        \data_from_adc[2]_104 , \data_from_adc[1]_81 , 
        \data_from_adc[1]_82 , \data_from_adc[1]_83 , 
        \data_from_adc[1]_84 , \data_from_adc[1]_85 , 
        \data_from_adc[4]_128 , \data_from_adc[3]_105 , 
        \data_from_adc[3]_106 , \data_from_adc[3]_107 , 
        \data_from_adc[3]_108 , \data_from_adc[3]_109 , 
        \data_from_adc[3]_110 , \data_from_adc[3]_111 , 
        \data_from_adc[3]_112 , \data_from_adc[3]_113 , 
        \data_from_adc[3]_114 , \data_from_adc[3]_115 , 
        \data_from_adc[3]_116 , \data_from_adc[2]_93 , 
        \data_from_adc[2]_94 , \data_from_adc[5]_137 , 
        \data_from_adc[5]_138 , \data_from_adc[5]_139 , 
        \data_from_adc[5]_140 , \data_from_adc[4]_117 , 
        \data_from_adc[4]_118 , \data_from_adc[4]_119 , 
        \data_from_adc[4]_120 , \data_from_adc[4]_121 , 
        \data_from_adc[4]_122 , \data_from_adc[4]_123 , 
        \data_from_adc[4]_124 , \data_from_adc[4]_125 , 
        \data_from_adc[4]_126 , \data_from_adc[4]_127 , temp1_15, 
        temp1_16, temp1_17, \cnt_frame[0]_net_1 , N_76_i_0, 
        \cnt_frame[1]_net_1 , N_74_i_0, \cnt_frame[2]_net_1 , N_72_i_0, 
        \cnt_frame[3]_net_1 , \cnt_frame_0_0[3]_net_1 , 
        \data_from_adc[5]_129 , \data_from_adc[5]_130 , 
        \data_from_adc[5]_131 , \data_from_adc[5]_132 , 
        \data_from_adc[5]_133 , \data_from_adc[5]_134 , 
        \data_from_adc[5]_135 , \data_from_adc[5]_136 , temp2_32, 
        temp2_33, temp1_2, temp1_3, temp1_4, temp1_5, temp1_6, temp1_7, 
        temp1_8, temp1_9, temp1_10, temp1_11, temp1_12, temp1_13, 
        temp1_14, temp2_18, temp2_19, temp2_20, temp2_21, temp2_22, 
        temp2_23, temp2_24, temp2_25, temp2_26, temp2_27, temp2_28, 
        temp2_29, temp2_30, temp2_31, clk_dac1_2_net_1, N_37_i_0, 
        N_35_i_0, SENSE_CS_1_4_iv_i_0, state15, N_13_i_0, freq15, 
        \un1_data_from_adc[2]_2_i_0 , \dac_count_1[7] , 
        clk_dac14_net_1, \dac_count_1[6] , \dac_count_3[5]_net_1 , 
        \dac_count_3[4]_net_1 , \dac_count_3[3]_net_1 , 
        \dac_count_3[2]_net_1 , \dac_count_3[1]_net_1 , cnt_freq6, 
        \cnt_freq[1]_net_1 , \cnt_freq_s[1] , \cnt_freq[2]_net_1 , 
        \cnt_freq_s[2] , \cnt_freq[3]_net_1 , \cnt_freq_s[3] , 
        \cnt_freq[4]_net_1 , \cnt_freq_s[4] , \cnt_freq[5]_net_1 , 
        \cnt_freq_s[5] , \cnt_freq[6]_net_1 , \cnt_freq_s[6] , 
        \cnt_freq[7]_net_1 , \cnt_freq_s[7] , \cnt_freq[8]_net_1 , 
        \cnt_freq_s[8] , \cnt_freq[9]_net_1 , \cnt_freq_s[9] , 
        \cnt_freq[10]_net_1 , \cnt_freq_s[10] , \cnt_freq[11]_net_1 , 
        \cnt_freq_s[11] , \cnt_freq[12]_net_1 , \cnt_freq_s[12] , 
        \cnt_freq[13]_net_1 , \cnt_freq_s[13] , \cnt_freq[14]_net_1 , 
        \cnt_freq_s[14] , \cnt_freq[15]_net_1 , \cnt_freq_s[15] , 
        \cnt_freq[16]_net_1 , \cnt_freq_s[16] , \cnt_freq[17]_net_1 , 
        \cnt_freq_s[17] , \cnt_freq[18]_net_1 , \cnt_freq_s[18] , 
        \cnt_freq[19]_net_1 , \cnt_freq_s[19] , \cnt_freq[20]_net_1 , 
        \cnt_freq_s[20] , \cnt_freq[21]_net_1 , \cnt_freq_s[21] , 
        \cnt_freq[22]_net_1 , \cnt_freq_s[22] , \cnt_freq[23]_net_1 , 
        \cnt_freq_s[23] , \cnt_freq[24]_net_1 , \cnt_freq_s[24] , 
        \cnt_freq[25]_net_1 , \cnt_freq_s[25] , \cnt_freq[26]_net_1 , 
        \cnt_freq_s[26] , \cnt_freq[27]_net_1 , \cnt_freq_s[27] , 
        \cnt_freq[28]_net_1 , \cnt_freq_s[28] , \cnt_freq[29]_net_1 , 
        \cnt_freq_s[29] , \cnt_freq[30]_net_1 , \cnt_freq_s[30] , 
        \cnt_freq[31]_net_1 , \cnt_freq_s[31]_net_1 , \cnt_s[0] , cnte, 
        \cnt[1]_net_1 , \cnt_s[1] , \cnt[2]_net_1 , \cnt_s[2] , 
        \cnt[3]_net_1 , \cnt_s[3] , \cnt[4]_net_1 , \cnt_s[4] , 
        \cnt[5]_net_1 , \cnt_s[5]_net_1 , \temp_count_s[0] , 
        \temp_count_s[1] , \temp_count_s[2] , \temp_count_s[3] , 
        \temp_count_s[4] , \temp_count_s[5] , \temp_count_s[6] , 
        \temp_count_s[7] , \temp_count_s[8] , \temp_count_s[9] , 
        \temp_count_s[10] , \temp_count_s[11] , \temp_count_s[12] , 
        \temp_count_s[13] , \temp_count_s[14] , \temp_count_s[15] , 
        \temp_count_s[16] , \temp_count_s[17] , \temp_count_s[18] , 
        \temp_count_s[19] , \temp_count_s[20] , \temp_count_s[21] , 
        \temp_count_s[22] , \temp_count_s[23] , \temp_count_s[24] , 
        \temp_count_s[25] , \temp_count_s[26] , \temp_count_s[27] , 
        \temp_count_s[28] , \temp_count_s[29] , \temp_count_s[30] , 
        \temp_count_s[31] , \fpga_count_s[1] , \fpga_count_s[2] , 
        \fpga_count_s[3] , \fpga_count_s[4] , \fpga_count_s[5] , 
        \fpga_count_s[6] , \fpga_count_s[7] , \fpga_count_s[8] , 
        \fpga_count_s[9] , \fpga_count_s[10] , \fpga_count_s[11] , 
        \fpga_count_s[12] , \fpga_count_s[13] , 
        \fpga_count_s[14]_net_1 , fpga_flags, N_109, 
        temp3_csn_RNO_net_1, un1_temp_state_7_or, 
        temp2_csn_RNO_0_net_1, un1_temp_state29_3_or, 
        temp1_csn_RNO_net_1, un1_temp_state_8_or, cnt_cry_cy, 
        un1_cnt_frame_0_sqmuxa_0_net_1, \cnt_cry[0]_net_1 , 
        \cnt_cry[1]_net_1 , \cnt_cry[2]_net_1 , \cnt_cry[3]_net_1 , 
        \cnt_cry[4]_net_1 , temp_count_lcry_cy, temp_count_net_1, 
        temp_count6_cry_31_RNIPJ5K1_Y, temp_count6, 
        \temp_count_cry[0] , \temp_count_cry[1] , \temp_count_cry[2] , 
        \temp_count_cry[3] , \temp_count_cry[4] , \temp_count_cry[5] , 
        \temp_count_cry[6] , \temp_count_cry[7] , \temp_count_cry[8] , 
        \temp_count_cry[9] , \temp_count_cry[10] , 
        \temp_count_cry[11] , \temp_count_cry[12] , 
        \temp_count_cry[13] , \temp_count_cry[14] , 
        \temp_count_cry[15] , \temp_count_cry[16] , 
        \temp_count_cry[17] , \temp_count_cry[18] , 
        \temp_count_cry[19] , \temp_count_cry[20] , 
        \temp_count_cry[21] , \temp_count_cry[22] , 
        \temp_count_cry[23] , \temp_count_cry[24] , 
        \temp_count_cry[25] , \temp_count_cry[26] , 
        \temp_count_cry[27] , \temp_count_cry[28] , 
        \temp_count_cry[29] , \temp_count_cry[30] , 
        dac_count_1_cry_0_net_1, dac_count_1_cry_0_Y, 
        dac_count_1_cry_1_net_1, \dac_count_1[2] , 
        dac_count_1_cry_2_net_1, \dac_count_1[3] , 
        dac_count_1_cry_3_net_1, \dac_count_1[4] , 
        dac_count_1_cry_4_net_1, \dac_count_1[5] , 
        dac_count_1_cry_5_net_1, un1_fr_adc_count_1_cry_1_net_1, 
        un1_fr_adc_count_1_cry_2_net_1, un1_fr_adc_count_1_cry_3_net_1, 
        un1_fr_adc_count_1_cry_4_net_1, un1_fr_adc_count_1_cry_5_net_1, 
        un1_fr_adc_count_1_cry_6_net_1, un1_fr_adc_count_1_cry_7_net_1, 
        un1_fr_adc_count_cry_1_net_1, un1_fr_adc_count_cry_2_net_1, 
        un1_fr_adc_count_cry_3_net_1, un1_fr_adc_count_cry_4_net_1, 
        un1_fr_adc_count_cry_5_net_1, un1_fr_adc_count_cry_6_net_1, 
        un1_fr_adc_count_cry_7_net_1, cnt_freq6_cry_7_net_1, 
        cnt_freq6_cry_8_net_1, cnt_freq6_cry_9_net_1, 
        cnt_freq6_cry_10_net_1, cnt_freq6_cry_11_net_1, 
        cnt_freq6_cry_12_net_1, cnt_freq6_cry_13_net_1, 
        cnt_freq6_cry_14_net_1, cnt_freq6_cry_15_net_1, 
        cnt_freq6_cry_16_net_1, cnt_freq6_cry_17_net_1, 
        cnt_freq6_cry_18_net_1, cnt_freq6_cry_19_net_1, 
        cnt_freq6_cry_20_net_1, cnt_freq6_cry_21_net_1, 
        cnt_freq6_cry_22_net_1, cnt_freq6_cry_23_net_1, 
        cnt_freq6_cry_24_net_1, cnt_freq6_cry_25_net_1, 
        cnt_freq6_cry_26_net_1, cnt_freq6_cry_27_net_1, 
        cnt_freq6_cry_28_net_1, cnt_freq6_cry_29_net_1, 
        cnt_freq6_cry_30_net_1, temp_count6_cry_7_net_1, 
        temp_count6_cry_8_net_1, temp_count6_cry_9_net_1, 
        temp_count6_cry_10_net_1, temp_count6_cry_11_net_1, 
        temp_count6_cry_12_net_1, temp_count6_cry_13_net_1, 
        temp_count6_cry_14_net_1, temp_count6_cry_15_net_1, 
        temp_count6_cry_16_net_1, temp_count6_cry_17_net_1, 
        temp_count6_cry_18_net_1, temp_count6_cry_19_net_1, 
        temp_count6_cry_20_net_1, temp_count6_cry_21_net_1, 
        temp_count6_cry_22_net_1, temp_count6_cry_23_net_1, 
        temp_count6_cry_24_net_1, temp_count6_cry_25_net_1, 
        temp_count6_cry_26_net_1, temp_count6_cry_27_net_1, 
        temp_count6_cry_28_net_1, temp_count6_cry_29_net_1, 
        temp_count6_cry_30_net_1, \fpga_flag4_0_data_tmp[0] , 
        \fpga_flag4_0_data_tmp[1] , \fpga_flag4_0_data_tmp[2] , 
        \fpga_flag4_0_data_tmp[3] , \fpga_flag4_0_data_tmp[4] , 
        \fpga_flag4_0_data_tmp[5] , \fpga_flag4_0_data_tmp[6] , 
        fpga_count_s_530_FCO, \fpga_count_cry[1]_net_1 , 
        \fpga_count_cry[2]_net_1 , \fpga_count_cry[3]_net_1 , 
        \fpga_count_cry[4]_net_1 , \fpga_count_cry[5]_net_1 , 
        \fpga_count_cry[6]_net_1 , \fpga_count_cry[7]_net_1 , 
        \fpga_count_cry[8]_net_1 , \fpga_count_cry[9]_net_1 , 
        \fpga_count_cry[10]_net_1 , \fpga_count_cry[11]_net_1 , 
        \fpga_count_cry[12]_net_1 , \fpga_count_cry[13]_net_1 , 
        cnt_freq_s_531_FCO, \cnt_freq_cry[1]_net_1 , 
        \cnt_freq_cry[2]_net_1 , \cnt_freq_cry[3]_net_1 , 
        \cnt_freq_cry[4]_net_1 , \cnt_freq_cry[5]_net_1 , 
        \cnt_freq_cry[6]_net_1 , \cnt_freq_cry[7]_net_1 , 
        \cnt_freq_cry[8]_net_1 , \cnt_freq_cry[9]_net_1 , 
        \cnt_freq_cry[10]_net_1 , \cnt_freq_cry[11]_net_1 , 
        \cnt_freq_cry[12]_net_1 , \cnt_freq_cry[13]_net_1 , 
        \cnt_freq_cry[14]_net_1 , \cnt_freq_cry[15]_net_1 , 
        \cnt_freq_cry[16]_net_1 , \cnt_freq_cry[17]_net_1 , 
        \cnt_freq_cry[18]_net_1 , \cnt_freq_cry[19]_net_1 , 
        \cnt_freq_cry[20]_net_1 , \cnt_freq_cry[21]_net_1 , 
        \cnt_freq_cry[22]_net_1 , \cnt_freq_cry[23]_net_1 , 
        \cnt_freq_cry[24]_net_1 , \cnt_freq_cry[25]_net_1 , 
        \cnt_freq_cry[26]_net_1 , \cnt_freq_cry[27]_net_1 , 
        \cnt_freq_cry[28]_net_1 , \cnt_freq_cry[29]_net_1 , 
        \cnt_freq_cry[30]_net_1 , N_10, m7_am, m7_bm, 
        \un1_data_from_adc[2]lt10 , \un1_data_from_adc[2]_2lt10 , 
        freq3lt11, data_m1_e_0_1, GPIO3_6_net_1, N_47, N_52, N_105, 
        N_2, N_170, N_73, N_51, freq3lt8, 
        \data_from_adc[0]_69_0_0_a2_1 , 
        \un1_data_from_adc[2]_1lto11_i_a2_7_net_1 , 
        \un1_data_from_adc[2]_1lto11_i_a2_6_net_1 , 
        \un1_data_from_adc[2]_1lto11_i_a2_5_net_1 , 
        \SENSE_DOUT_2_1_u_i_a3_3_0[1]_net_1 , freq3lto8_1_net_1, 
        \SENSE_DOUT_2_1_u_i_a3_0[1]_net_1 , 
        \cnt_frame_0_0_a3_0_1_0[3]_net_1 , GPIO3_9_net_1, 
        GPIO3_8_net_1, GPIO3_7_net_1, GPIO5_13_net_1, GPIO5_12_net_1, 
        GPIO5_11_net_1, GPIO5_10_net_1, 
        \data_from_adc[4]_0_sqmuxa_3_net_1 , un22_data_from_adc_net_1, 
        \data_from_adc[7]_0_sqmuxa_3_net_1 , 
        \data_from_adc[5]_0_sqmuxa_3_net_1 , 
        \data_from_adc[3]_0_sqmuxa_3_net_1 , 
        \data_from_adc[1]_0_sqmuxa_3_net_1 , N_48, 
        \data_from_adc[6]_0_sqmuxa_3_net_1 , SENSE_CS_1_1_sqmuxalt5, 
        un12_data_from_adc_net_1, un14_data_from_adc_net_1, 
        un13_data_from_adc_net_1, N_123, un18_data_from_adc_net_1, 
        \un1_data_from_adc[2]lto8_0_net_1 , _decfrac4, 
        un15_data_from_adc_net_1, un20_data_from_adc_net_1, 
        un21_data_from_adc_net_1, N_82, N_168, N_49, N_50, N_129, N_90, 
        N_183, \un1_data_from_adc[2]lt5 , GPIO5_14_net_1, 
        \data_from_adc[2]_0_sqmuxa_0_a2_3_RNO_net_1 , N_125, N_185, 
        N_714, \SENSE_DOUT_2_1_u_i_1[1]_net_1 , 
        \SENSE_DOUT_2_1_u_i_0[1]_net_1 , N_130, N_96;
    
    SLE \cnt[0]  (.D(\cnt_s[0] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(GPIO7_c));
    SLE \SENSE_DOUT_1[1]  (.D(N_37_i_0), .CLK(temp_sck_c_i_0), .EN(
        N_35_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(SENSE_DOUT_c[1]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[3]_114 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(N_185), .Y(
        \data_from_adc[8]_166 ));
    SLE \data_from_adc[1][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_91 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [10]));
    CFG3 #( .INIT(8'h41) )  \temp_count_data_RNO[2]  (.A(
        temp_count_data[4]), .B(temp_count_data[2]), .C(N_73), .Y(
        N_11_i_0));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[4]_128 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[7]_164 ));
    SLE fpga_flag (.D(fpga_flags), .CLK(BW_clk_c_i_0), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(fpga_flag_i), .SD(
        VCC_net_1), .LAT(GND_net_1), .Q(fpga_flag_net_1));
    SLE \temp_count_data[3]  (.D(N_9_i_0), .CLK(temp_sck_c), .EN(
        un1_temp_state28_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count_data[3]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(N_183), .C(N_96), .Y(
        \data_from_adc[2]_102 ));
    ARI1 #( .INIT(20'h555AA) )  dac_count_1_cry_3 (.A(dac_count[4]), 
        .B(fr_adc_count[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_1_cry_2_net_1), .S(\dac_count_1[4] ), .Y(), .FCO(
        dac_count_1_cry_3_net_1));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_21 (.A(freq_14), .B(
        \cnt_freq[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_20_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_21_net_1));
    SLE \temp_count[14]  (.D(\temp_count_s[14] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[14]));
    SLE \BW_out[13]  (.D(fpga_count[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[13]));
    ARI1 #( .INIT(20'h42200) )  \temp_state_RNIL54L[2]  (.A(VCC_net_1), 
        .B(\temp_state[1]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        GND_net_1), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        temp_count_lcry_cy));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNICB9I61[18]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[18]), .D(GND_net_1), .FCI(\temp_count_cry[17] ), .S(
        \temp_count_s[18] ), .Y(), .FCO(\temp_count_cry[18] ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_23 (.A(VCC_net_1), .B(
        \cnt_freq[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_22_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_23_net_1));
    SLE \data_from_adc[7][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_157 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [4]));
    CFG4 #( .INIT(16'h0800) )  temp3_34_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_50), .Y(temp3_34));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[12]  (.A(VCC_net_1), .B(
        \cnt_freq[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[11]_net_1 ), .S(\cnt_freq_s[12] ), .Y(), .FCO(
        \cnt_freq_cry[12]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \cnt_freq_RNO[0]  (.A(\cnt_freq[0]_net_1 ), 
        .Y(\cnt_freq_s[0] ));
    SLE \dac1_db[12]  (.D(dac1_db_8_6_236_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[12]));
    SLE \cnt_freq[11]  (.D(\cnt_freq_s[11] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[11]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_21 (.A(freq_14), .B(
        temp_count[21]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_20_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_21_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[11]  (.A(VCC_net_1), .B(
        \cnt_freq[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[10]_net_1 ), .S(\cnt_freq_s[11] ), .Y(), .FCO(
        \cnt_freq_cry[11]_net_1 ));
    SLE \data_from_adc[5][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_137 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [8]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(N_183), .C(N_96), .Y(
        \data_from_adc[2]_104 ));
    SLE \fpga_count[0]  (.D(\fpga_count_s[0] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[0]));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[1]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(\data_from_adc[1]_0_sqmuxa_3_net_1 ), 
        .Y(\data_from_adc[1]_87 ));
    SLE \temp3[1]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_35), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[1]));
    SLE \fpga_shift_2[7]  (.D(BW_out_c[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[7]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[2]  (.A(VCC_net_1), .B(
        \cnt_freq[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[1]_net_1 ), .S(\cnt_freq_s[2] ), .Y(), .FCO(
        \cnt_freq_cry[2]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_2_276_i_m2 (.A(dds_cos[3]), .B(
        sdv_count[1]), .C(dds_sin[3]), .Y(dac1_db_8_2_276_i_m2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[18]  (.A(VCC_net_1), .B(
        \cnt_freq[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[17]_net_1 ), .S(\cnt_freq_s[18] ), .Y(), .FCO(
        \cnt_freq_cry[18]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(N_125), .Y(
        \data_from_adc[0]_71 ));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[6]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(\data_from_adc[6]_0_sqmuxa_3_net_1 ), 
        .Y(\data_from_adc[6]_147 ));
    CFG4 #( .INIT(16'h0001) )  \SENSE_DOUT_2_1_u_i_a3_2[1]  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(N_125));
    SLE \data_from_adc[7][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_162 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [9]));
    CFG1 #( .INIT(2'h1) )  clk_dac1_2_RNO (.A(sdv_count[1]), .Y(
        \sdv_count_i_0[1] ));
    SLE \BW_out[2]  (.D(fpga_count[2]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[2]));
    SLE \data_from_adc[2][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_93 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [0]));
    CFG4 #( .INIT(16'h0051) )  freq9 (.A(\data_from_adc[2] [11]), .B(
        \data_from_adc[2] [10]), .C(\un1_data_from_adc[2]lt10 ), .D(
        freq3), .Y(freq9_net_1));
    SLE \BW_out[8]  (.D(fpga_count[8]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[8]));
    SLE \BW_out[0]  (.D(fpga_count[0]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[0]));
    CFG4 #( .INIT(16'h0010) )  temp2_18_0_0_a2 (.A(temp_count_data[4]), 
        .B(\temp_state[0]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(N_48));
    SLE \cnt_freq[27]  (.D(\cnt_freq_s[27] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[27]_net_1 ));
    SLE \data_from_adc[4][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_123 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [6]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6US111[15]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[15]), .D(GND_net_1), .FCI(\temp_count_cry[14] ), .S(
        \temp_count_s[15] ), .Y(), .FCO(\temp_count_cry[15] ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6O6JH1[24]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[24]), .D(GND_net_1), .FCI(\temp_count_cry[23] ), .S(
        \temp_count_s[24] ), .Y(), .FCO(\temp_count_cry[24] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[3]_115 ));
    CFG4 #( .INIT(16'h0C09) )  \cnt_frame_RNO[2]  (.A(N_105), .B(
        \cnt_frame[2]_net_1 ), .C(N_129), .D(N_90), .Y(N_72_i_0));
    SLE \temp_count[30]  (.D(\temp_count_s[30] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[30]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[3]  (.A(VCC_net_1), .B(
        \cnt_freq[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[2]_net_1 ), .S(\cnt_freq_s[3] ), .Y(), .FCO(
        \cnt_freq_cry[3]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_4_256_i_m2 (.A(dds_cos[5]), .B(
        sdv_count[1]), .C(dds_sin[5]), .Y(dac1_db_8_4_256_i_m2_net_1));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[7]_RNO[8]  (.A(N_82), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(N_168), .Y(
        \data_from_adc[7]_161 ));
    SLE \BW_out[10]  (.D(fpga_count[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[10]));
    SLE \temp2[13]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_31), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[13]));
    SLE \freq[17]  (.D(freq3_i_0), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_10));
    CFG4 #( .INIT(16'h0200) )  temp1_6_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_49), .Y(temp1_6));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[4]  (.A(VCC_net_1), .B(
        un1_cnt_frame_0_sqmuxa_0_net_1), .C(\cnt[4]_net_1 ), .D(
        GND_net_1), .FCI(\cnt_cry[3]_net_1 ), .S(\cnt_s[4] ), .Y(), 
        .FCO(\cnt_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_12 (.A(freq_2), .B(
        temp_count[12]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_11_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_12_net_1));
    SLE \data_from_adc[2][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_98 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [5]));
    SLE \fpga_shift_2[13]  (.D(BW_out_c[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[13]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_11 (.A(freq_1), .B(
        \cnt_freq[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_10_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_11_net_1));
    SLE \temp_count[2]  (.D(\temp_count_s[2] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[2]));
    SLE \temp_count[27]  (.D(\temp_count_s[27] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[27]));
    SLE \dac_count[1]  (.D(\dac_count_3[1]_net_1 ), .CLK(BW_clk_c), 
        .EN(clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[1]));
    SLE \data_from_adc[6][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_151 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [10]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(N_125), .C(N_96), .Y(
        \data_from_adc[0]_76 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_13 (.A(freq_6), .B(
        \cnt_freq[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_12_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_13_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI5I897[2]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[2]), .D(
        GND_net_1), .FCI(\temp_count_cry[1] ), .S(\temp_count_s[2] ), 
        .Y(), .FCO(\temp_count_cry[2] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_fr_adc_count_cry_7 (.A(VCC_net_1), 
        .B(dac_count[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_fr_adc_count_cry_6_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_cry_7_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[20]  (.A(VCC_net_1), .B(
        \cnt_freq[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[19]_net_1 ), .S(\cnt_freq_s[20] ), .Y(), .FCO(
        \cnt_freq_cry[20]_net_1 ));
    SLE \cnt_freq[5]  (.D(\cnt_freq_s[5] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[5]_net_1 ));
    SLE \temp3[11]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_45), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[11]));
    CFG4 #( .INIT(16'h2000) )  temp3_45_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_50), .D(N_47), .Y(temp3_45));
    SLE temp1_csn (.D(\temp_state[0]_net_1 ), .CLK(temp_sck_c), .EN(
        temp1_csn_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_449_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(temp1_csn_c));
    SLE \data_from_adc[6][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_152 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [11]));
    SLE \data_from_adc[3][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_107 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [2]));
    CFG4 #( .INIT(16'h0100) )  temp3_46_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_50), .Y(temp3_46));
    SLE \data_from_adc[7][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_161 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [8]));
    CFG4 #( .INIT(16'h0010) )  \SENSE_DOUT_2_1_u_i_a3_0[1]  (.A(
        \cnt_frame[1]_net_1 ), .B(\cnt[1]_net_1 ), .C(
        \cnt_frame[0]_net_1 ), .D(GPIO7_c), .Y(N_123));
    SLE \cnt_freq[17]  (.D(\cnt_freq_s[17] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[17]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \un1_data_from_adc[2]lto4  (.A(
        \data_from_adc[2] [2]), .B(\data_from_adc[2] [4]), .C(
        \data_from_adc[2] [3]), .Y(\un1_data_from_adc[2]lt5 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIG7URN[10]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[10]), .D(GND_net_1), .FCI(\temp_count_cry[9] ), .S(
        \temp_count_s[10] ), .Y(), .FCO(\temp_count_cry[10] ));
    SLE \fpga_shift_2[4]  (.D(BW_out_c[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[4]));
    CFG2 #( .INIT(4'h2) )  \dac_count_3[2]  (.A(\dac_count_1[2] ), .B(
        un1_fr_adc_count_cry_7_net_1), .Y(\dac_count_3[2]_net_1 ));
    SLE \dac_count[2]  (.D(\dac_count_3[2]_net_1 ), .CLK(BW_clk_c), 
        .EN(clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[2]));
    CFG2 #( .INIT(4'h1) )  temp_count_data_n0_i_a3 (.A(
        temp_count_data[4]), .B(temp_count_data[0]), .Y(N_33));
    CFG3 #( .INIT(8'h02) )  \SENSE_DOUT_2_1_u_i_a3_3_0[1]  (.A(
        \cnt_frame[2]_net_1 ), .B(\cnt_frame[1]_net_1 ), .C(
        \cnt_frame[0]_net_1 ), .Y(\SENSE_DOUT_2_1_u_i_a3_3_0[1]_net_1 )
        );
    CFG4 #( .INIT(16'h6996) )  GPIO5_10 (.A(GPS1_I0_c), .B(GPIO9_c), 
        .C(GPIO6_c), .D(GPIO4_c), .Y(GPIO5_10_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[14]  (.A(VCC_net_1), .B(
        \cnt_freq[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[13]_net_1 ), .S(\cnt_freq_s[14] ), .Y(), .FCO(
        \cnt_freq_cry[14]_net_1 ));
    SLE \dac_count[5]  (.D(\dac_count_3[5]_net_1 ), .CLK(BW_clk_c), 
        .EN(clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[5]));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_6_236_i_m2 (.A(dds_cos[7]), .B(
        sdv_count[1]), .C(dds_sin[7]), .Y(dac1_db_8_6_236_i_m2_net_1));
    SLE \temp2[2]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_20), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[2]));
    CFG4 #( .INIT(16'hFCFE) )  \data_from_adc[2]_0_sqmuxa_0_a2_3  (.A(
        \data_from_adc[0]_69_0_0_a2_1 ), .B(N_168), .C(
        \data_from_adc[2]_0_sqmuxa_0_a2_3_RNO_net_1 ), .D(N_82), .Y(
        N_96));
    SLE \data_from_adc[2][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_97 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [4]));
    SLE \data_from_adc[1][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_83 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [2]));
    SLE \data_from_adc[0][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_72 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [3]));
    CFG1 #( .INIT(2'h1) )  \fpga_count_RNO[0]  (.A(fpga_count[0]), .Y(
        \fpga_count_s[0] ));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[3]  (.A(VCC_net_1), .B(
        un1_cnt_frame_0_sqmuxa_0_net_1), .C(\cnt[3]_net_1 ), .D(
        GND_net_1), .FCI(\cnt_cry[2]_net_1 ), .S(\cnt_s[3] ), .Y(), 
        .FCO(\cnt_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI0Q2GB[4]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[4]), .D(
        GND_net_1), .FCI(\temp_count_cry[3] ), .S(\temp_count_s[4] ), 
        .Y(), .FCO(\temp_count_cry[4] ));
    SLE \fpga_count[3]  (.D(\fpga_count_s[3] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[3]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[13]  (.A(VCC_net_1), 
        .B(fpga_count[13]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[12]_net_1 ), .S(\fpga_count_s[13] ), .Y(), 
        .FCO(\fpga_count_cry[13]_net_1 ));
    SLE \temp1[15]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_17), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[15]));
    SLE \fpga_count[5]  (.D(\fpga_count_s[5] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[5]));
    SLE \temp1[2]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_4), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[2]));
    SLE \temp3[12]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_46), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[12]));
    ARI1 #( .INIT(20'h65500) )  un1_fr_adc_count_1_cry_7 (.A(VCC_net_1)
        , .B(dac_count[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_fr_adc_count_1_cry_6_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_1_cry_7_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[1]  (.A(VCC_net_1), .B(
        \cnt_freq[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq_s_531_FCO), .S(\cnt_freq_s[1] ), .Y(), .FCO(
        \cnt_freq_cry[1]_net_1 ));
    SLE \cnt[3]  (.D(\cnt_s[3] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[3]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[5]  (.A(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .B(_decfrac4), .C(N_96), 
        .Y(\data_from_adc[4]_122 ));
    SLE \fpga_shift_2[12]  (.D(BW_out_c[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[12]));
    SLE \temp2[14]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_32), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[14]));
    SLE \data_from_adc[4][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_127 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [10]));
    CFG4 #( .INIT(16'h4000) )  temp2_25_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_48), .D(N_47), .Y(temp2_25));
    CFG3 #( .INIT(8'hFE) )  SENSE_DOUT61_i_o2 (.A(\cnt[2]_net_1 ), .B(
        \cnt[1]_net_1 ), .C(GPIO7_c), .Y(N_82));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[5]_133 ));
    SLE \data_from_adc[2][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_102 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [9]));
    SLE SENSE_CS_1 (.D(SENSE_CS_1_4_iv_i_0), .CLK(temp_sck_c_i_0), .EN(
        state15), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(SENSE_CS_1_c));
    ARI1 #( .INIT(20'h49900) )  fpga_flag4_0_I_45 (.A(VCC_net_1), .B(
        fpga_shift_2[14]), .C(\fpga_data_receive[14]_net_1 ), .D(
        GND_net_1), .FCI(\fpga_flag4_0_data_tmp[6] ), .S(), .Y(), .FCO(
        fpga_flags));
    CFG4 #( .INIT(16'h0400) )  temp2_26_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_48), .Y(temp2_26));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_10 (.A(freq_0), .B(
        temp_count[10]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_9_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_10_net_1));
    CFG3 #( .INIT(8'hFB) )  \cnt_frame_0_i_o2[0]  (.A(\state[1]_net_1 )
        , .B(\state[0]_net_1 ), .C(\cnt_frame[3]_net_1 ), .Y(N_90));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_1_cry_2 (.A(
        dac_count[2]), .B(fr_adc_count[2]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_fr_adc_count_1_cry_1_net_1), .S(), .Y(), 
        .FCO(un1_fr_adc_count_1_cry_2_net_1));
    CFG4 #( .INIT(16'h0040) )  \temp_count_data_RNO[4]  (.A(
        temp_count_data[4]), .B(temp_count_data[3]), .C(
        temp_count_data[2]), .D(N_73), .Y(N_7_i_0));
    CFG4 #( .INIT(16'h3310) )  \un1_data_from_adc[2]lto9  (.A(
        \data_from_adc[2] [5]), .B(\data_from_adc[2] [9]), .C(
        \un1_data_from_adc[2]lt5 ), .D(
        \un1_data_from_adc[2]lto8_0_net_1 ), .Y(
        \un1_data_from_adc[2]lt10 ));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_27 (.A(
        \fpga_data_receive[7]_net_1 ), .B(fpga_shift_2[6]), .C(
        fpga_shift_2[7]), .D(\fpga_data_receive[6]_net_1 ), .FCI(
        \fpga_flag4_0_data_tmp[2] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[3] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[3]_106 ));
    SLE \data_from_adc[3][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_115 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [10]));
    CFG3 #( .INIT(8'h4E) )  \temp_state_7_2_0_.m7_bm  (.A(
        temp_count_data[4]), .B(\temp_state[0]_net_1 ), .C(
        \temp_state[1]_net_1 ), .Y(m7_bm));
    CFG1 #( .INIT(2'h1) )  temp2_csn_RNO (.A(\temp_state[1]_net_1 ), 
        .Y(\temp_state_i_0[1] ));
    SLE \cnt_freq[20]  (.D(\cnt_freq_s[20] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[20]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI7THTD1[22]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[22]), .D(GND_net_1), .FCI(\temp_count_cry[21] ), .S(
        \temp_count_s[22] ), .Y(), .FCO(\temp_count_cry[22] ));
    SLE \temp3[6]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_40), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[6]));
    SLE \fpga_data_receive[13]  (.D(BW_c[13]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[13]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[7]_0_sqmuxa_3  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ));
    SLE \temp2[10]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_28), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[10]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIFVFJD[5]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[5]), .D(
        GND_net_1), .FCI(\temp_count_cry[4] ), .S(\temp_count_s[5] ), 
        .Y(), .FCO(\temp_count_cry[5] ));
    SLE \fpga_count[8]  (.D(\fpga_count_s[8] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[8]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(N_183), .Y(
        \data_from_adc[2]_94 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(N_183), .C(N_96), .Y(
        \data_from_adc[2]_103 ));
    SLE \temp3[0]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_34), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[0]));
    CFG4 #( .INIT(16'h8000) )  \un1_data_from_adc[2]_1lto11_i_a2_5  (
        .A(\data_from_adc[2] [1]), .B(\data_from_adc[2] [0]), .C(
        \data_from_adc[2] [6]), .D(\data_from_adc[2] [5]), .Y(
        \un1_data_from_adc[2]_1lto11_i_a2_5_net_1 ));
    CFG4 #( .INIT(16'h6996) )  GPIO3_9 (.A(adc_d0_c[11]), .B(
        adc_d0_c[10]), .C(adc_d0_c[9]), .D(adc_d0_c[8]), .Y(
        GPIO3_9_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNICGNMP[11]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[11]), .D(GND_net_1), .FCI(\temp_count_cry[10] ), .S(
        \temp_count_s[11] ), .Y(), .FCO(\temp_count_cry[11] ));
    CFG3 #( .INIT(8'h01) )  \state_5_i_i_a3[0]  (.A(\state[0]_net_1 ), 
        .B(GPIO11_c), .C(\state[1]_net_1 ), .Y(N_129));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_23 (.A(VCC_net_1), .B(
        temp_count[23]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_22_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_23_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[5]  (.A(_decfrac4), 
        .B(N_96), .C(N_185), .Y(\data_from_adc[8]_170 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(N_125), .C(N_96), .Y(
        \data_from_adc[0]_79 ));
    SLE \cnt_freq[24]  (.D(\cnt_freq_s[24] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[24]_net_1 ));
    SLE \cnt_freq[22]  (.D(\cnt_freq_s[22] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[22]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIGDAQH[7]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[7]), .D(
        GND_net_1), .FCI(\temp_count_cry[6] ), .S(\temp_count_s[7] ), 
        .Y(), .FCO(\temp_count_cry[7] ));
    CFG2 #( .INIT(4'h2) )  \dac_count_3[5]  (.A(\dac_count_1[5] ), .B(
        un1_fr_adc_count_cry_7_net_1), .Y(\dac_count_3[5]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[7]_155 ));
    SLE \data_from_adc[2][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_101 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [8]));
    SLE \temp2[5]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_23), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[5]));
    SLE \data_from_adc[4][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_118 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [1]));
    SLE \temp2[7]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_25), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[7]));
    SLE \cnt_frame[3]  (.D(\cnt_frame_0_0[3]_net_1 ), .CLK(
        temp_sck_c_i_0), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\cnt_frame[3]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[5]_138 ));
    SLE \BW_out[6]  (.D(fpga_count[6]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[6]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNO[31]  (.A(VCC_net_1), 
        .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[31]), .D(
        GND_net_1), .FCI(\temp_count_cry[30] ), .S(\temp_count_s[31] ), 
        .Y(), .FCO());
    SLE \data_from_adc[5][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_132 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [3]));
    CFG2 #( .INIT(4'h4) )  state15_0_a2 (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(state15));
    SLE \data_from_adc[4][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_124 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [7]));
    SLE \temp1[7]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_9), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[7]));
    SLE \dac_count[7]  (.D(\dac_count_1[7] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[7]));
    SLE \cnt_freq[10]  (.D(\cnt_freq_s[10] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[10]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIILLC9[3]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[3]), .D(
        GND_net_1), .FCI(\temp_count_cry[2] ), .S(\temp_count_s[3] ), 
        .Y(), .FCO(\temp_count_cry[3] ));
    SLE \fpga_data_receive[7]  (.D(BW_c[7]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[7]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[4]_RNO[8]  (.A(N_82), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(N_168), .Y(
        \data_from_adc[4]_125 ));
    SLE \data_from_adc[0][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_75 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [6]));
    SLE \temp_count[23]  (.D(\temp_count_s[23] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[23]));
    SLE \cnt_freq[9]  (.D(\cnt_freq_s[9] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[9]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_29 (.A(VCC_net_1), .B(
        \cnt_freq[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_28_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_29_net_1));
    SLE \temp_count[17]  (.D(\temp_count_s[17] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[17]));
    SLE \cnt_freq[14]  (.D(\cnt_freq_s[14] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[14]_net_1 ));
    SLE \cnt_freq[12]  (.D(\cnt_freq_s[12] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[12]_net_1 ));
    SLE \cnt_freq[26]  (.D(\cnt_freq_s[26] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[26]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[1]_85 ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_14 (.A(VCC_net_1), .B(
        temp_count[14]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_13_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_14_net_1));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_30 (.A(VCC_net_1), .B(
        temp_count[30]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_29_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_30_net_1));
    CFG4 #( .INIT(16'h1000) )  \data_from_adc[3]_0_sqmuxa_3  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[15]  (.A(VCC_net_1), .B(
        \cnt_freq[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[14]_net_1 ), .S(\cnt_freq_s[15] ), .Y(), .FCO(
        \cnt_freq_cry[15]_net_1 ));
    SLE \fpga_shift_2[11]  (.D(BW_out_c[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[11]));
    CFG4 #( .INIT(16'h0004) )  \data_from_adc[4]_0_sqmuxa_3  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[7]_160 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[6]_145 ));
    ARI1 #( .INIT(20'h6AA00) )  temp_count6_cry_19 (.A(VCC_net_1), .B(
        temp_count[19]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_18_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_19_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIC8M3N1[27]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[27]), .D(GND_net_1), .FCI(\temp_count_cry[26] ), .S(
        \temp_count_s[27] ), .Y(), .FCO(\temp_count_cry[27] ));
    SLE \sdv_count[1]  (.D(\sdv_count_1[1] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(sdv_count[1]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNILV41M[9]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[9]), .D(
        GND_net_1), .FCI(\temp_count_cry[8] ), .S(\temp_count_s[9] ), 
        .Y(), .FCO(\temp_count_cry[9] ));
    SLE \freq[21]  (.D(\fr_adc_count_5_i_0[2] ), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_14));
    SLE \temp2[8]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_26), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[8]));
    CFG4 #( .INIT(16'h0080) )  un13_data_from_adc (.A(\cnt[3]_net_1 ), 
        .B(\cnt[2]_net_1 ), .C(\cnt[1]_net_1 ), .D(GPIO7_c), .Y(
        un13_data_from_adc_net_1));
    SLE \fpga_shift_2[3]  (.D(BW_out_c[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[3]));
    SLE \fpga_shift_2[1]  (.D(BW_out_c[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[1]));
    SLE \data_from_adc[2][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_104 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [11]));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[8]_RNO[8]  (.A(N_82), .B(
        N_185), .C(N_168), .Y(\data_from_adc[8]_173 ));
    CFG4 #( .INIT(16'h3C20) )  temp2_csn_RNO_1 (.A(temp_count_data[4]), 
        .B(\temp_state[0]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(un1_temp_state29_3_or));
    SLE \data_from_adc[7][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_156 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [3]));
    CFG3 #( .INIT(8'hA3) )  \temp_state_7_2_0_.N_11_i  (.A(
        \temp_state[0]_net_1 ), .B(N_10), .C(\temp_state[2]_net_1 ), 
        .Y(N_11_i_0_0));
    CFG3 #( .INIT(8'h40) )  \cnt_frame_0_0_a3_0_1_0[3]  (.A(
        \state[1]_net_1 ), .B(\state[0]_net_1 ), .C(
        \cnt_frame[2]_net_1 ), .Y(\cnt_frame_0_0_a3_0_1_0[3]_net_1 ));
    SLE \cnt_freq[16]  (.D(\cnt_freq_s[16] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[16]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  dac_count_1_cry_5 (.A(VCC_net_1), .B(
        dac_count[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_1_cry_4_net_1), .S(\dac_count_1[6] ), .Y(), .FCO(
        dac_count_1_cry_5_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[17]  (.A(VCC_net_1), .B(
        \cnt_freq[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[16]_net_1 ), .S(\cnt_freq_s[17] ), .Y(), .FCO(
        \cnt_freq_cry[17]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  GPIO5_12 (.A(GPS_I0_c), .B(GPS2_Q1_c), 
        .C(GPS2_Q0_c), .D(GPS2_LD_c), .Y(GPIO5_12_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[1]_90 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(N_125), .Y(
        \data_from_adc[0]_72 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_17 (.A(freq_10), .B(
        temp_count[17]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_16_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_17_net_1));
    dds dds_w (.dds_sin({dds_sin[7], dds_sin[6], dds_sin[5], 
        dds_sin[4], dds_sin[3], dds_sin[2], dds_sin[1], dds_sin[0]}), 
        .dds_cos({dds_cos[7], dds_cos[6], dds_cos[5], dds_cos[4], 
        dds_cos[3], dds_cos[2], dds_cos[1], dds_cos[0]}), .dac_count({
        dac_count[7], dac_count[6], dac_count[5], dac_count[4], 
        dac_count[3], dac_count[2], dac_count[1]}), .BW_clk_c(BW_clk_c)
        );
    ARI1 #( .INIT(20'h6AA00) )  cnt_freq6_cry_19 (.A(VCC_net_1), .B(
        \cnt_freq[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_18_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_19_net_1));
    CFG2 #( .INIT(4'h2) )  _decfrac4_0_a2 (.A(\cnt[1]_net_1 ), .B(
        \cnt[2]_net_1 ), .Y(N_170));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_28 (.A(VCC_net_1), .B(
        \cnt_freq[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_27_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_28_net_1));
    SLE \cnt_freq[25]  (.D(\cnt_freq_s[25] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[25]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  temp1_8_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_49), .Y(temp1_8));
    CFG4 #( .INIT(16'h8000) )  temp1_3_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_49), .Y(temp1_3));
    SLE \cnt_frame[2]  (.D(N_72_i_0), .CLK(temp_sck_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_frame[2]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[6]_150 ));
    SLE \temp_count[9]  (.D(\temp_count_s[9] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[9]));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_8 (.A(freq_1), .B(
        temp_count[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_7_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_8_net_1));
    SLE \data_from_adc[5][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_135 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [6]));
    SLE \cnt_freq[31]  (.D(\cnt_freq_s[31]_net_1 ), .CLK(temp_sck_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        cnt_freq6), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \cnt_freq[31]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  temp3_35_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_50), .Y(temp3_35));
    CFG4 #( .INIT(16'h8000) )  temp3_36_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_50), .Y(temp3_36));
    SLE \dac_count[6]  (.D(\dac_count_1[6] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[6]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_9 (.A(freq_2), .B(
        \cnt_freq[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_8_net_1), .S(), .Y(), .FCO(cnt_freq6_cry_9_net_1)
        );
    CFG2 #( .INIT(4'h8) )  _decfrac4_0_a3 (.A(N_170), .B(GPIO7_c), .Y(
        _decfrac4));
    SLE \data_from_adc[8][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_175 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [10]));
    CFG2 #( .INIT(4'h6) )  \sdv_count_RNO[1]  (.A(sdv_count[1]), .B(
        sdv_count[0]), .Y(\sdv_count_1[1] ));
    SLE \dac1_db[5]  (.D(dac1_db_8_306_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[5]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[26]  (.A(VCC_net_1), .B(
        \cnt_freq[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[25]_net_1 ), .S(\cnt_freq_s[26] ), .Y(), .FCO(
        \cnt_freq_cry[26]_net_1 ));
    CFG4 #( .INIT(16'hFC54) )  \SENSE_DOUT_2_1_u_i_a3_0_1[1]  (.A(
        \cnt_frame[2]_net_1 ), .B(\cnt_frame[1]_net_1 ), .C(
        \cnt_frame[0]_net_1 ), .D(GPIO7_c), .Y(
        \SENSE_DOUT_2_1_u_i_a3_0[1]_net_1 ));
    SLE \temp_count[6]  (.D(\temp_count_s[6] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[6]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI7CMS21[16]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[16]), .D(GND_net_1), .FCI(\temp_count_cry[15] ), .S(
        \temp_count_s[16] ), .Y(), .FCO(\temp_count_cry[16] ));
    ARI1 #( .INIT(20'h4AA00) )  dac_count_1_s_6 (.A(VCC_net_1), .B(
        dac_count[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_1_cry_5_net_1), .S(\dac_count_1[7] ), .Y(), .FCO());
    CFG1 #( .INIT(2'h1) )  temp_state26_0_a3_RNIBC45 (.A(temp_state26), 
        .Y(N_449_i));
    SLE \data_from_adc[8][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_165 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [0]));
    ARI1 #( .INIT(20'h4AAA2) )  \temp_count_RNIEEE23[0]  (.A(
        temp_count6), .B(temp_count[0]), .C(\temp_state[1]_net_1 ), .D(
        \temp_state[2]_net_1 ), .FCI(temp_count_net_1), .S(
        \temp_count_s[0] ), .Y(), .FCO(\temp_count_cry[0] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[1]_92 ));
    SLE \cnt_freq[15]  (.D(\cnt_freq_s[15] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[15]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[1]_91 ));
    ARI1 #( .INIT(20'h555AA) )  dac_count_1_cry_1 (.A(dac_count[2]), 
        .B(fr_adc_count[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_1_cry_0_net_1), .S(\dac_count_1[2] ), .Y(), .FCO(
        dac_count_1_cry_1_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9NR8L1[26]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[26]), .D(GND_net_1), .FCI(\temp_count_cry[25] ), .S(
        \temp_count_s[26] ), .Y(), .FCO(\temp_count_cry[26] ));
    SLE \temp1[13]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_15), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[13]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[4]_119 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[19]  (.A(VCC_net_1), .B(
        \cnt_freq[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[18]_net_1 ), .S(\cnt_freq_s[19] ), .Y(), .FCO(
        \cnt_freq_cry[19]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \data_from_adc[0]_RNO[0]  (.A(N_125), .B(
        \data_from_adc[0]_69_0_0_a2_1 ), .C(N_82), .Y(
        \data_from_adc[0]_69 ));
    SLE \dac1_db[11]  (.D(dac1_db_8_5_246_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[11]));
    SLE \BW_out[9]  (.D(fpga_count[9]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[9]));
    SLE \fpga_data_receive[8]  (.D(BW_c[8]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[8]_net_1 ));
    SLE \cnt_freq[0]  (.D(\cnt_freq_s[0] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[0]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[5]  (.A(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .B(_decfrac4), .C(N_96), 
        .Y(\data_from_adc[3]_110 ));
    SLE \data_from_adc[8][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_170 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [5]));
    SLE \temp1[6]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_8), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[6]));
    SLE \data_from_adc[4][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_119 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [2]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_18 (.A(freq_11), .B(
        \cnt_freq[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_17_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_18_net_1));
    SLE \data_from_adc[0][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_70 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [1]));
    SLE \temp3[9]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_43), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[9]));
    CFG2 #( .INIT(4'hB) )  \fr_adc_count_5_0_a2_i[2]  (.A(freq3), .B(
        \un1_data_from_adc[2]_2 ), .Y(\fr_adc_count_5_i_0[2] ));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_306_i_m2 (.A(dds_cos[0]), .B(
        sdv_count[1]), .C(dds_sin[0]), .Y(dac1_db_8_306_i_m2_net_1));
    SLE \temp_count[13]  (.D(\temp_count_s[13] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[13]));
    SLE \data_from_adc[2][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_96 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [3]));
    SLE \data_from_adc[7][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_159 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [6]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[5]  (.A(_decfrac4), 
        .B(N_96), .C(N_183), .Y(\data_from_adc[2]_98 ));
    SLE \fpga_shift_2[0]  (.D(BW_out_c[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[0]));
    SLE \data_from_adc[0][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_76 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [7]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[5]_130 ));
    SLE \data_from_adc[5][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_140 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [11]));
    ARI1 #( .INIT(20'h4AA00) )  un1_fr_adc_count_cry_6 (.A(VCC_net_1), 
        .B(dac_count[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_fr_adc_count_cry_5_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_cry_6_net_1));
    CFG4 #( .INIT(16'h0010) )  \data_from_adc[2]_0_sqmuxa_0_a2_0  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(N_183));
    SLE \temp2[9]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_27), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[9]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[6]_151 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_s[31]  (.A(VCC_net_1), .B(
        \cnt_freq[31]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[30]_net_1 ), .S(\cnt_freq_s[31]_net_1 ), .Y(), 
        .FCO());
    SLE \data_from_adc[3][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_116 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [11]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_27 (.A(VCC_net_1), .B(
        \cnt_freq[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_26_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_27_net_1));
    SLE \fpga_count[1]  (.D(\fpga_count_s[1] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[1]));
    SLE \temp1[5]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_7), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[5]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[4]_124 ));
    SLE \temp_state[1]  (.D(N_11_i_0_0), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\temp_state[1]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(N_185), .Y(
        \data_from_adc[8]_167 ));
    SLE \fpga_shift_2[10]  (.D(BW_out_c[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[10]));
    SLE \cnt_freq[28]  (.D(\cnt_freq_s[28] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[28]_net_1 ));
    SLE \fpga_data_receive[4]  (.D(BW_c[4]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[4]_net_1 ));
    SLE \data_from_adc[8][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_169 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [4]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI75ACT[13]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[13]), .D(GND_net_1), .FCI(\temp_count_cry[12] ), .S(
        \temp_count_s[13] ), .Y(), .FCO(\temp_count_cry[13] ));
    SLE \BW_out[1]  (.D(fpga_count[1]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[1]));
    SLE \temp_count[21]  (.D(\temp_count_s[21] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[21]));
    CFG2 #( .INIT(4'h4) )  temp2_27_0_0_a2 (.A(temp_count_data[0]), .B(
        temp_count_data[1]), .Y(N_52));
    CFG3 #( .INIT(8'h7F) )  
        \un1_data_from_adc[2]_1lto11_i_a2_5_RNI4DVM  (.A(
        \un1_data_from_adc[2]_1lto11_i_a2_6_net_1 ), .B(
        \un1_data_from_adc[2]_1lto11_i_a2_7_net_1 ), .C(
        \un1_data_from_adc[2]_1lto11_i_a2_5_net_1 ), .Y(
        \un1_data_from_adc[2]_1_i_i_0 ));
    SLE \temp_count[22]  (.D(\temp_count_s[22] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[22]));
    CFG4 #( .INIT(16'h0800) )  \data_from_adc[0]_RNO[6]  (.A(N_168), 
        .B(N_125), .C(GPIO7_c), .D(N_170), .Y(\data_from_adc[0]_75 ));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[2]  (.A(VCC_net_1), .B(
        un1_cnt_frame_0_sqmuxa_0_net_1), .C(\cnt[2]_net_1 ), .D(
        GND_net_1), .FCI(\cnt_cry[1]_net_1 ), .S(\cnt_s[2] ), .Y(), 
        .FCO(\cnt_cry[2]_net_1 ));
    CFG4 #( .INIT(16'hFEEE) )  SENSE_CS_1_1_sqmuxalto3 (.A(
        \cnt[3]_net_1 ), .B(\cnt[2]_net_1 ), .C(\cnt[1]_net_1 ), .D(
        GPIO7_c), .Y(SENSE_CS_1_1_sqmuxalt5));
    SLE \temp1[14]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_16), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[14]));
    SLE \freq[22]  (.D(\un1_data_from_adc[2]_i_0 ), .CLK(temp_sck_c), 
        .EN(\un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_15));
    SLE \data_from_adc[8][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_174 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [9]));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[3]_RNO[8]  (.A(N_82), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(N_168), .Y(
        \data_from_adc[3]_113 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(N_185), .C(N_96), .Y(
        \data_from_adc[8]_172 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[7]_156 ));
    SLE \data_from_adc[5][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_130 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [1]));
    SLE \cnt_freq[18]  (.D(\cnt_freq_s[18] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[18]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_fr_adc_count_1_cry_6 (.A(VCC_net_1)
        , .B(dac_count[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_fr_adc_count_1_cry_5_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_1_cry_6_net_1));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[2]_RNO[8]  (.A(N_82), .B(
        N_183), .C(N_168), .Y(\data_from_adc[2]_101 ));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_9 (.A(
        \fpga_data_receive[13]_net_1 ), .B(fpga_shift_2[12]), .C(
        fpga_shift_2[13]), .D(\fpga_data_receive[12]_net_1 ), .FCI(
        \fpga_flag4_0_data_tmp[5] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[6] ));
    SLE \data_from_adc[6][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_141 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [0]));
    SLE \data_from_adc[5][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_136 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [7]));
    CFG3 #( .INIT(8'h7F) )  \un1_data_from_adc[2]lto8_0  (.A(
        \data_from_adc[2] [8]), .B(\data_from_adc[2] [7]), .C(
        \data_from_adc[2] [6]), .Y(\un1_data_from_adc[2]lto8_0_net_1 ));
    SLE \temp1[10]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_12), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[10]));
    SLE \fr_adc_count[2]  (.D(\fr_adc_count_5[2] ), .CLK(temp_sck_c), 
        .EN(\un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fr_adc_count[2]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_17 (.A(freq_10), .B(
        \cnt_freq[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_16_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_17_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .Y(\data_from_adc[1]_82 )
        );
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_1_286_i_m2 (.A(dds_cos[2]), .B(
        sdv_count[1]), .C(dds_sin[2]), .Y(dac1_db_8_1_286_i_m2_net_1));
    CFG4 #( .INIT(16'hFFF7) )  freq3lto8 (.A(\data_from_adc[2] [7]), 
        .B(\data_from_adc[2] [8]), .C(freq3lto8_1_net_1), .D(freq3lt8), 
        .Y(freq3lt11));
    SLE \data_from_adc[2][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_99 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [6]));
    SLE \temp_count_data[0]  (.D(N_33), .CLK(temp_sck_c), .EN(
        un1_temp_state28_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count_data[0]));
    CFG4 #( .INIT(16'h2000) )  temp1_13_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_49), .D(N_47), .Y(temp1_13));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[6]_142 ));
    SLE \fr_adc_count[1]  (.D(\fr_adc_count_5[1] ), .CLK(temp_sck_c), 
        .EN(\un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fr_adc_count[1]));
    SLE \data_from_adc[6][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_146 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [5]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9RFN41[17]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[17]), .D(GND_net_1), .FCI(\temp_count_cry[16] ), .S(
        \temp_count_s[17] ), .Y(), .FCO(\temp_count_cry[17] ));
    CFG4 #( .INIT(16'h8CC0) )  temp3_csn_RNO_0 (.A(temp_count_data[4]), 
        .B(\temp_state[0]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(un1_temp_state_7_or));
    CFG4 #( .INIT(16'h0800) )  temp1_2_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_49), .Y(temp1_2));
    SLE \data_from_adc[8][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_173 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [8]));
    CFG4 #( .INIT(16'hFFAE) )  freq9_i_0 (.A(\data_from_adc[2] [11]), 
        .B(\data_from_adc[2] [10]), .C(\un1_data_from_adc[2]lt10 ), .D(
        freq3), .Y(freq9_i_0_net_1));
    CFG4 #( .INIT(16'h151F) )  \temp_state_7_2_0_.m9  (.A(
        \temp_state[0]_net_1 ), .B(temp_count6), .C(
        \temp_state[1]_net_1 ), .D(temp_count_data[4]), .Y(N_10));
    SLE \temp_state[0]  (.D(\temp_state_7[0] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\temp_state[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un12_data_from_adc (.A(\cnt[3]_net_1 ), 
        .B(\cnt[2]_net_1 ), .C(\cnt[1]_net_1 ), .D(GPIO7_c), .Y(
        un12_data_from_adc_net_1));
    CFG2 #( .INIT(4'h1) )  temp_count_data_n1_i_a2 (.A(
        temp_count_data[0]), .B(temp_count_data[1]), .Y(N_47));
    SLE \cnt_freq[30]  (.D(\cnt_freq_s[30] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[30]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  un14_data_from_adc (.A(\cnt[3]_net_1 ), 
        .B(\cnt[2]_net_1 ), .C(\cnt[1]_net_1 ), .D(GPIO7_c), .Y(
        un14_data_from_adc_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[23]  (.A(VCC_net_1), .B(
        \cnt_freq[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[22]_net_1 ), .S(\cnt_freq_s[23] ), .Y(), .FCO(
        \cnt_freq_cry[23]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \dac_count_3[1]  (.A(
        un1_fr_adc_count_cry_7_net_1), .B(dac_count_1_cry_0_Y), .Y(
        \dac_count_3[1]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_9 (.A(freq_2), .B(
        temp_count[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_8_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_9_net_1));
    CFG4 #( .INIT(16'h0100) )  \data_from_adc[1]_0_sqmuxa_3  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ));
    CFG2 #( .INIT(4'hE) )  \fr_adc_count_5_0[1]  (.A(freq15), .B(freq3)
        , .Y(\fr_adc_count_5[1] ));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_1 (.A(
        \fpga_data_receive[1]_net_1 ), .B(fpga_shift_2[0]), .C(
        fpga_shift_2[1]), .D(\fpga_data_receive[0]_net_1 ), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(\fpga_flag4_0_data_tmp[0] ));
    SLE \temp_count[3]  (.D(\temp_count_s[3] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[3]));
    SLE \fpga_data_receive[2]  (.D(BW_c[2]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[8]  (.A(VCC_net_1), .B(
        fpga_count[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[7]_net_1 ), .S(\fpga_count_s[8] ), .Y(), .FCO(
        \fpga_count_cry[8]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[7]_RNO[0]  (.A(N_82), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(
        \data_from_adc[0]_69_0_0_a2_1 ), .Y(\data_from_adc[7]_153 ));
    SLE \data_from_adc[7][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_154 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [1]));
    SLE \data_from_adc[7][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_163 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [10]));
    SLE \dac1_db[10]  (.D(dac1_db_8_4_256_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[10]));
    SLE temp3_csn (.D(N_109), .CLK(temp_sck_c), .EN(
        temp3_csn_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_449_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(temp3_csn_c));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[8]  (.A(VCC_net_1), .B(
        \cnt_freq[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[7]_net_1 ), .S(\cnt_freq_s[8] ), .Y(), .FCO(
        \cnt_freq_cry[8]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_7 (.A(freq_0), .B(
        \cnt_freq[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(cnt_freq6_cry_7_net_1));
    SLE \data_from_adc[7][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_160 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [7]));
    SLE \fpga_data_receive[11]  (.D(BW_c[11]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[11]_net_1 ));
    SLE \data_from_adc[6][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_145 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [4]));
    SLE \data_from_adc[0][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_71 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [2]));
    SLE \freq[13]  (.D(freq15), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_6));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_26 (.A(VCC_net_1), .B(
        temp_count[26]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_25_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_26_net_1));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_20 (.A(freq_13), .B(
        \cnt_freq[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_19_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_20_net_1));
    SLE \fpga_count[4]  (.D(\fpga_count_s[4] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[4]));
    ARI1 #( .INIT(20'h555AA) )  dac_count_1_cry_0 (.A(dac_count[1]), 
        .B(fr_adc_count[1]), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(dac_count_1_cry_0_Y), .FCO(
        dac_count_1_cry_0_net_1));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_24 (.A(VCC_net_1), .B(
        \cnt_freq[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_23_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_24_net_1));
    SLE \fpga_shift_2[8]  (.D(BW_out_c[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[8]));
    CFG4 #( .INIT(16'hFEFF) )  freq3lto11_i (.A(\data_from_adc[2] [9]), 
        .B(\data_from_adc[2] [11]), .C(\data_from_adc[2] [10]), .D(
        freq3lt11), .Y(freq3_i_0));
    CFG4 #( .INIT(16'h0004) )  temp1_2_0_0_a2 (.A(temp_count_data[4]), 
        .B(\temp_state[0]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(N_49));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_28 (.A(VCC_net_1), .B(
        temp_count[28]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_27_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_28_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[3]_116 ));
    SLE \data_from_adc[6][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_150 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [9]));
    CFG2 #( .INIT(4'h2) )  temp2_24_0_0_a2 (.A(temp_count_data[0]), .B(
        temp_count_data[1]), .Y(N_51));
    SLE \temp3[7]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_41), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[7]));
    SLE \temp_count[11]  (.D(\temp_count_s[11] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[11]));
    CFG3 #( .INIT(8'h02) )  un15_data_from_adc (.A(\cnt[2]_net_1 ), .B(
        \cnt[1]_net_1 ), .C(GPIO7_c), .Y(un15_data_from_adc_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[5]_140 ));
    SLE \dac1_db[13]  (.D(dac1_db_0_sqmuxa_net_1), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[13]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_22 (.A(freq_15), .B(
        \cnt_freq[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_21_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_22_net_1));
    SLE \temp_count[12]  (.D(\temp_count_s[12] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[12]));
    SLE \fpga_data_receive[1]  (.D(BW_c[1]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \un1_data_from_adc[2]_1lto11_i_a2_6  (
        .A(\data_from_adc[2] [9]), .B(\data_from_adc[2] [4]), .C(
        \data_from_adc[2] [10]), .D(\data_from_adc[2] [11]), .Y(
        \un1_data_from_adc[2]_1lto11_i_a2_6_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6ACOF1[23]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[23]), .D(GND_net_1), .FCI(\temp_count_cry[22] ), .S(
        \temp_count_s[23] ), .Y(), .FCO(\temp_count_cry[23] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[3]_107 ));
    SLE \fpga_count[6]  (.D(\fpga_count_s[6] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[6]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[5]  (.A(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .B(_decfrac4), .C(N_96), 
        .Y(\data_from_adc[5]_134 ));
    SLE \temp3[15]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_49), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[15]));
    CFG4 #( .INIT(16'h4000) )  temp1_11_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_49), .Y(temp1_11));
    CFG2 #( .INIT(4'h4) )  dac1_db_0_sqmuxa (.A(
        un1_fr_adc_count_1_cry_7_net_1), .B(sdv_count[1]), .Y(
        dac1_db_0_sqmuxa_net_1));
    SLE \temp1[0]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_2), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[0]));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_cry_4 (.A(
        dac_count[4]), .B(fr_adc_count[2]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_fr_adc_count_cry_3_net_1), .S(), .Y(), 
        .FCO(un1_fr_adc_count_cry_4_net_1));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[7]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(\data_from_adc[7]_0_sqmuxa_3_net_1 ), 
        .Y(\data_from_adc[7]_159 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(N_183), .Y(
        \data_from_adc[2]_95 ));
    SLE \fr_adc_count[5]  (.D(\un1_data_from_adc[2]_2_i_0 ), .CLK(
        temp_sck_c), .EN(\un1_data_from_adc[2]_1_i_i_0 ), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(freq_2));
    SLE \temp_count[25]  (.D(\temp_count_s[25] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[25]));
    SLE \temp2[11]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_29), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[11]));
    CFG4 #( .INIT(16'h4000) )  temp3_34_0_0_a2 (.A(temp_count_data[4]), 
        .B(\temp_state[0]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(N_50));
    SLE \data_from_adc[3][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_105 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [0]));
    SLE \BW_out[5]  (.D(fpga_count[5]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[5]));
    SLE \fpga_data_receive[0]  (.D(BW_c[0]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[0]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \data_from_adc[2]_0_sqmuxa_0_a2_3_RNO_0  (
        .A(\cnt[4]_net_1 ), .B(\cnt[5]_net_1 ), .Y(data_m1_e_0_1));
    SLE \data_from_adc[6][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_149 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [8]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[4]_120 ));
    SLE \state[1]  (.D(N_40_i_0), .CLK(temp_sck_c_i_0), .EN(
        un1_state15_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state[1]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_10 (.A(freq_0), .B(
        \cnt_freq[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_9_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_10_net_1));
    SLE \dac_count[4]  (.D(\dac_count_3[4]_net_1 ), .CLK(BW_clk_c), 
        .EN(clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[4]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_14 (.A(VCC_net_1), .B(
        \cnt_freq[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_13_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_14_net_1));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_15 (.A(freq_0), .B(
        temp_count[15]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_14_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_15_net_1));
    SLE \temp_count[26]  (.D(\temp_count_s[26] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[26]));
    SLE \data_from_adc[5][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_131 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [2]));
    CFG4 #( .INIT(16'h6996) )  GPIO3_8 (.A(adc_d0_c[7]), .B(
        adc_d0_c[6]), .C(adc_d0_c[5]), .D(adc_d0_c[4]), .Y(
        GPIO3_8_net_1));
    SLE \data_from_adc[2][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_94 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [1]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6H37V[14]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[14]), .D(GND_net_1), .FCI(\temp_count_cry[13] ), .S(
        \temp_count_s[14] ), .Y(), .FCO(\temp_count_cry[14] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[3]_112 ));
    CFG3 #( .INIT(8'h10) )  \data_from_adc[2]_0_sqmuxa_0_a2_1  (.A(
        \cnt[5]_net_1 ), .B(\cnt[4]_net_1 ), .C(\cnt[3]_net_1 ), .Y(
        N_168));
    SLE \data_from_adc[1][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_81 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [0]));
    SLE \data_from_adc[3][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_110 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [5]));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[1]  (.A(VCC_net_1), .B(
        un1_cnt_frame_0_sqmuxa_0_net_1), .C(\cnt[1]_net_1 ), .D(
        GND_net_1), .FCI(\cnt_cry[0]_net_1 ), .S(\cnt_s[1] ), .Y(), 
        .FCO(\cnt_cry[1]_net_1 ));
    SLE \data_from_adc[2][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_100 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [7]));
    SLE \dac1_db[9]  (.D(dac1_db_8_3_266_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[9]));
    CFG4 #( .INIT(16'h3733) )  \un1_data_from_adc[2]_2lto11  (.A(
        \data_from_adc[2] [9]), .B(\data_from_adc[2] [11]), .C(
        \data_from_adc[2] [10]), .D(\un1_data_from_adc[2]_2lt10 ), .Y(
        \un1_data_from_adc[2]_2 ));
    CFG3 #( .INIT(8'h10) )  un18_data_from_adc (.A(\cnt[2]_net_1 ), .B(
        \cnt[1]_net_1 ), .C(GPIO7_c), .Y(un18_data_from_adc_net_1));
    CFG4 #( .INIT(16'hAE00) )  \fr_adc_count_5_0_a2[1]  (.A(
        \data_from_adc[2] [11]), .B(\data_from_adc[2] [10]), .C(
        \un1_data_from_adc[2]lt10 ), .D(\un1_data_from_adc[2]_2 ), .Y(
        freq15));
    SLE \data_from_adc[8][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_176 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [11]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(N_125), .C(N_96), .Y(
        \data_from_adc[0]_73 ));
    CFG4 #( .INIT(16'h4000) )  temp3_43_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_50), .Y(temp3_43));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(N_183), .C(N_96), .Y(
        \data_from_adc[2]_100 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[5]  (.A(VCC_net_1), .B(
        fpga_count[5]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[4]_net_1 ), .S(\fpga_count_s[5] ), .Y(), .FCO(
        \fpga_count_cry[5]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_12 (.A(freq_2), .B(
        \cnt_freq[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_11_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_12_net_1));
    SLE \temp_count[1]  (.D(\temp_count_s[1] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[1]));
    SLE \temp2[12]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_30), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[12]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[11]  (.A(VCC_net_1), 
        .B(fpga_count[11]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[10]_net_1 ), .S(\fpga_count_s[11] ), .Y(), 
        .FCO(\fpga_count_cry[11]_net_1 ));
    SLE \cnt[4]  (.D(\cnt_s[4] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[4]_net_1 ));
    ARI1 #( .INIT(20'h4EF00) )  temp_count6_cry_31_RNIPJ5K1 (.A(
        VCC_net_1), .B(temp_count6), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .FCI(temp_count_lcry_cy), .S(), .Y(
        temp_count6_cry_31_RNIPJ5K1_Y), .FCO(temp_count_net_1));
    SLE \freq[7]  (.D(freq9_net_1), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_0));
    CFG3 #( .INIT(8'h41) )  \cnt_frame_RNO[0]  (.A(N_129), .B(
        \cnt_frame[0]_net_1 ), .C(N_90), .Y(N_76_i_0));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[4]_127 ));
    ARI1 #( .INIT(20'h4AA00) )  cnt_freq_s_531 (.A(VCC_net_1), .B(
        \cnt_freq[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(cnt_freq_s_531_FCO));
    SLE \data_from_adc[1][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_86 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [5]));
    SLE \cnt_freq[2]  (.D(\cnt_freq_s[2] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[2]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_31 (.A(VCC_net_1), .B(
        \cnt_freq[31]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_30_net_1), .S(), .Y(), .FCO(cnt_freq6));
    CFG1 #( .INIT(2'h1) )  fpga_flag_RNO (.A(fpga_flag_net_1), .Y(
        fpga_flag_i));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(N_185), .Y(
        \data_from_adc[8]_168 ));
    SLE \cnt[5]  (.D(\cnt_s[5]_net_1 ), .CLK(temp_sck_c_i_0), .EN(cnte)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[5]_net_1 ));
    SLE \fpga_count[9]  (.D(\fpga_count_s[9] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[9]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIC6T7A1[20]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[20]), .D(GND_net_1), .FCI(\temp_count_cry[19] ), .S(
        \temp_count_s[20] ), .Y(), .FCO(\temp_count_cry[20] ));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[5]_RNO[8]  (.A(N_82), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(N_168), .Y(
        \data_from_adc[5]_137 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[10]  (.A(VCC_net_1), .B(
        \cnt_freq[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[9]_net_1 ), .S(\cnt_freq_s[10] ), .Y(), .FCO(
        \cnt_freq_cry[10]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_11 (.A(freq_1), .B(
        temp_count[11]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_10_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_11_net_1));
    CFG4 #( .INIT(16'hEE6E) )  SENSE_CS_1_4_iv_i (.A(\cnt[4]_net_1 ), 
        .B(\cnt[5]_net_1 ), .C(SENSE_CS_1_1_sqmuxalt5), .D(
        SENSE_CS_1_c), .Y(SENSE_CS_1_4_iv_i_0));
    SLE \data_from_adc[8][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_168 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [3]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[5]  (.A(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .B(_decfrac4), .C(N_96), 
        .Y(\data_from_adc[1]_86 ));
    SLE \data_from_adc[3][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_109 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [4]));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[4]_RNO[0]  (.A(N_82), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(
        \data_from_adc[0]_69_0_0_a2_1 ), .Y(\data_from_adc[4]_117 ));
    CFG4 #( .INIT(16'hFEF2) )  \SENSE_DOUT_2_1_0[1]  (.A(
        \cnt_frame[2]_net_1 ), .B(\cnt[2]_net_1 ), .C(GPIO7_c), .D(
        \cnt[1]_net_1 ), .Y(N_714));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9HN2C1[21]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[21]), .D(GND_net_1), .FCI(\temp_count_cry[20] ), .S(
        \temp_count_s[21] ), .Y(), .FCO(\temp_count_cry[21] ));
    CFG3 #( .INIT(8'h74) )  \temp_state_7_2_0_.m13  (.A(
        \temp_state[1]_net_1 ), .B(N_2), .C(\temp_state[2]_net_1 ), .Y(
        \temp_state_7[2] ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_22 (.A(freq_15), .B(
        temp_count[22]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_21_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_22_net_1));
    CFG4 #( .INIT(16'hF1F0) )  \un1_data_from_adc[2]_2lto8  (.A(
        \data_from_adc[2] [4]), .B(\data_from_adc[2] [5]), .C(
        \un1_data_from_adc[2]lto8_0_net_1 ), .D(freq3lt8), .Y(
        \un1_data_from_adc[2]_2lt10 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[5]  (.A(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .B(_decfrac4), .C(N_96), 
        .Y(\data_from_adc[6]_146 ));
    CFG1 #( .INIT(2'h1) )  \temp_state_RNI91IA[0]  (.A(
        \temp_state[0]_net_1 ), .Y(\temp_state_i_0[0] ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_26 (.A(VCC_net_1), .B(
        \cnt_freq[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_25_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_26_net_1));
    SLE \freq[20]  (.D(freq15_i_0), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_13));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[9]  (.A(VCC_net_1), .B(
        \cnt_freq[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[8]_net_1 ), .S(\cnt_freq_s[9] ), .Y(), .FCO(
        \cnt_freq_cry[9]_net_1 ));
    CFG4 #( .INIT(16'h51FF) )  \fr_adc_count_5_0_a2_i[1]  (.A(
        \data_from_adc[2] [11]), .B(\data_from_adc[2] [10]), .C(
        \un1_data_from_adc[2]lt10 ), .D(\un1_data_from_adc[2]_2 ), .Y(
        freq15_i_0));
    SLE \temp3[8]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_42), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[8]));
    SLE \data_from_adc[7][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_155 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [2]));
    CFG4 #( .INIT(16'h2000) )  temp2_23_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_48), .Y(temp2_23));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[22]  (.A(VCC_net_1), .B(
        \cnt_freq[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[21]_net_1 ), .S(\cnt_freq_s[22] ), .Y(), .FCO(
        \cnt_freq_cry[22]_net_1 ));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_33 (.A(
        \fpga_data_receive[5]_net_1 ), .B(fpga_shift_2[4]), .C(
        fpga_shift_2[5]), .D(\fpga_data_receive[4]_net_1 ), .FCI(
        \fpga_flag4_0_data_tmp[1] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[2] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(N_125), .C(N_96), .Y(
        \data_from_adc[0]_78 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[21]  (.A(VCC_net_1), .B(
        \cnt_freq[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[20]_net_1 ), .S(\cnt_freq_s[21] ), .Y(), .FCO(
        \cnt_freq_cry[21]_net_1 ));
    SLE \data_from_adc[3][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_114 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [9]));
    SLE \data_from_adc[1][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_85 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [4]));
    SLE \fpga_data_receive[6]  (.D(BW_c[6]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[6]_net_1 ));
    CFG2 #( .INIT(4'h8) )  clk_dac2_RNIJBB8 (.A(GPIO10_c), .B(clk_dac2)
        , .Y(dac2_clk_c));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[28]  (.A(VCC_net_1), .B(
        \cnt_freq[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[27]_net_1 ), .S(\cnt_freq_s[28] ), .Y(), .FCO(
        \cnt_freq_cry[28]_net_1 ));
    SLE \temp_count[20]  (.D(\temp_count_s[20] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[20]));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_15 (.A(
        \fpga_data_receive[11]_net_1 ), .B(fpga_shift_2[10]), .C(
        fpga_shift_2[11]), .D(\fpga_data_receive[10]_net_1 ), .FCI(
        \fpga_flag4_0_data_tmp[4] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[5] ));
    CFG4 #( .INIT(16'h6996) )  GPIO5_14 (.A(osc_vcc_c), .B(
        GPIO5_10_net_1), .C(ANTF_n2_c), .D(ANTF_n1_c), .Y(
        GPIO5_14_net_1));
    CFG4 #( .INIT(16'h8000) )  temp1_5_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_49), .D(N_47), .Y(temp1_5));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIV5TMF[6]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[6]), .D(
        GND_net_1), .FCI(\temp_count_cry[5] ), .S(\temp_count_s[6] ), 
        .Y(), .FCO(\temp_count_cry[6] ));
    CFG4 #( .INIT(16'hFF26) )  \state_RNIND411[0]  (.A(
        \state[1]_net_1 ), .B(\state[0]_net_1 ), .C(
        \cnt_frame[3]_net_1 ), .D(un1_cnt_frame_0_sqmuxa_0_net_1), .Y(
        cnte));
    SLE \temp1[9]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_11), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[9]));
    CFG3 #( .INIT(8'h08) )  \data_from_adc[8]_RNO[0]  (.A(N_185), .B(
        \data_from_adc[0]_69_0_0_a2_1 ), .C(N_82), .Y(
        \data_from_adc[8]_165 ));
    SLE \data_from_adc[1][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_90 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [9]));
    CFG2 #( .INIT(4'h7) )  un1_state15_0 (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(un1_state15_0_net_1));
    CFG4 #( .INIT(16'h3222) )  clk_dac1_2 (.A(\sdv_count_i_0[1] ), .B(
        clk_dac14_net_1), .C(dac1_clk_c), .D(sdv_count[1]), .Y(
        clk_dac1_2_net_1));
    CFG4 #( .INIT(16'h4000) )  temp1_12_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_49), .Y(temp1_12));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[5]_139 ));
    SLE \temp_count[8]  (.D(\temp_count_s[8] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[8]));
    CFG3 #( .INIT(8'hF2) )  \freq_RNO[22]  (.A(\data_from_adc[2] [10]), 
        .B(\un1_data_from_adc[2]lt10 ), .C(\data_from_adc[2] [11]), .Y(
        \un1_data_from_adc[2]_i_0 ));
    CFG2 #( .INIT(4'h1) )  clk_dac14 (.A(sdv_count[1]), .B(
        sdv_count[0]), .Y(clk_dac14_net_1));
    CFG4 #( .INIT(16'h4000) )  temp3_41_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_50), .D(N_47), .Y(temp3_41));
    SLE \fpga_count[13]  (.D(\fpga_count_s[13] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[13]));
    SLE \data_from_adc[0][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_80 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [11]));
    SLE \temp_count[15]  (.D(\temp_count_s[15] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[15]));
    SLE \temp2[1]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_19), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[1]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[2]  (.A(VCC_net_1), .B(
        fpga_count[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[1]_net_1 ), .S(\fpga_count_s[2] ), .Y(), .FCO(
        \fpga_count_cry[2]_net_1 ));
    SLE \sdv_count[0]  (.D(\sdv_count_i_0[0] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(sdv_count[0]));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[4]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(\data_from_adc[4]_0_sqmuxa_3_net_1 ), 
        .Y(\data_from_adc[4]_123 ));
    CFG4 #( .INIT(16'h0400) )  temp1_10_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_49), .Y(temp1_10));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[30]  (.A(VCC_net_1), .B(
        \cnt_freq[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[29]_net_1 ), .S(\cnt_freq_s[30] ), .Y(), .FCO(
        \cnt_freq_cry[30]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_31 (.A(VCC_net_1), .B(
        temp_count[31]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_30_net_1), .S(), .Y(), .FCO(temp_count6));
    SLE \data_from_adc[3][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_113 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [8]));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[1]_RNO[8]  (.A(N_82), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(N_168), .Y(
        \data_from_adc[1]_89 ));
    CFG4 #( .INIT(16'h1000) )  temp1_17_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_49), .D(N_47), .Y(temp1_17));
    SLE \temp1[4]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_6), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[4]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_16 (.A(freq_1), .B(
        \cnt_freq[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_15_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_16_net_1));
    CFG2 #( .INIT(4'hE) )  temp3_csn_RNO (.A(temp_state26), .B(
        un1_temp_state_7_or), .Y(temp3_csn_RNO_net_1));
    CFG2 #( .INIT(4'h7) )  \SENSE_DOUT_2_1_u_i_o2_3[1]  (.A(
        \cnt_frame[0]_net_1 ), .B(\cnt_frame[1]_net_1 ), .Y(N_105));
    CFG3 #( .INIT(8'h04) )  \cnt_RNIKLML[4]  (.A(\cnt[5]_net_1 ), .B(
        \cnt[4]_net_1 ), .C(\cnt[3]_net_1 ), .Y(
        \data_from_adc[0]_69_0_0_a2_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_20 (.A(freq_13), .B(
        temp_count[20]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_19_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_20_net_1));
    SLE \temp2[3]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_21), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[3]));
    CFG2 #( .INIT(4'hE) )  \state_5_i_i[0]  (.A(N_130), .B(N_129), .Y(
        N_42));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[6]_RNO[8]  (.A(N_82), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(N_168), .Y(
        \data_from_adc[6]_149 ));
    CFG2 #( .INIT(4'h2) )  \dac_count_3[3]  (.A(\dac_count_1[3] ), .B(
        un1_fr_adc_count_cry_7_net_1), .Y(\dac_count_3[3]_net_1 ));
    SLE \temp1[8]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_10), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[8]));
    SLE \temp_count[16]  (.D(\temp_count_s[16] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[16]));
    SLE \data_from_adc[8][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_171 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [6]));
    CFG2 #( .INIT(4'hE) )  temp2_csn_RNO_0 (.A(temp_state26), .B(
        un1_temp_state29_3_or), .Y(temp2_csn_RNO_0_net_1));
    CFG3 #( .INIT(8'h92) )  un1_temp_state28_0 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[1]_net_1 ), .C(
        \temp_state[0]_net_1 ), .Y(un1_temp_state28_0_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIPFR55[1]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[1]), .D(
        GND_net_1), .FCI(\temp_count_cry[0] ), .S(\temp_count_s[1] ), 
        .Y(), .FCO(\temp_count_cry[1] ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_7 (.A(freq_0), .B(
        temp_count[7]), .C(GND_net_1), .D(GND_net_1), .FCI(GND_net_1), 
        .S(), .Y(), .FCO(temp_count6_cry_7_net_1));
    SLE \data_from_adc[1][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_89 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [8]));
    SLE \BW_out[14]  (.D(fpga_count[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[14]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[24]  (.A(VCC_net_1), .B(
        \cnt_freq[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[23]_net_1 ), .S(\cnt_freq_s[24] ), .Y(), .FCO(
        \cnt_freq_cry[24]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(N_185), .C(N_96), .Y(
        \data_from_adc[8]_176 ));
    SLE \state[0]  (.D(N_42), .CLK(temp_sck_c_i_0), .EN(
        un1_state15_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state[0]_net_1 ));
    SLE \dac1_db[8]  (.D(dac1_db_8_2_276_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[8]));
    SLE \fpga_data_receive[9]  (.D(BW_c[9]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[9]_net_1 ));
    SLE \data_from_adc[6][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_144 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [3]));
    SLE \data_from_adc[2][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_95 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [2]));
    CFG2 #( .INIT(4'h8) )  \temp_state_7_2_0_.m1  (.A(
        \temp_state[0]_net_1 ), .B(temp_count_data[4]), .Y(N_2));
    CFG4 #( .INIT(16'h8000) )  temp2_21_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_48), .D(N_47), .Y(temp2_21));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[7]_157 ));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[8]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(N_185), .Y(\data_from_adc[8]_171 ));
    CFG4 #( .INIT(16'h1000) )  temp3_48_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_50), .Y(temp3_48));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[5]_131 ));
    CFG4 #( .INIT(16'hF8F0) )  \SENSE_DOUT_2_1_u_i_0[1]  (.A(N_105), 
        .B(N_170), .C(N_123), .D(\SENSE_DOUT_2_1_u_i_a3_0[1]_net_1 ), 
        .Y(\SENSE_DOUT_2_1_u_i_0[1]_net_1 ));
    CFG2 #( .INIT(4'h9) )  GPIO16_RNO (.A(cnt_freq6), .B(GPIO16_c), .Y(
        N_13_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[1]  (.A(VCC_net_1), .B(
        fpga_count[1]), .C(GND_net_1), .D(GND_net_1), .FCI(
        fpga_count_s_530_FCO), .S(\fpga_count_s[1] ), .Y(), .FCO(
        \fpga_count_cry[1]_net_1 ));
    SLE \cnt_freq[23]  (.D(\cnt_freq_s[23] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[23]_net_1 ));
    CFG3 #( .INIT(8'h04) )  un21_data_from_adc (.A(\cnt[3]_net_1 ), .B(
        \cnt[2]_net_1 ), .C(GPIO7_c), .Y(un21_data_from_adc_net_1));
    SLE \temp3[13]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_47), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[13]));
    CFG2 #( .INIT(4'h4) )  SENSE_CS_1_RNIM4KA (.A(SENSE_CS_1_c), .B(
        temp_sck_c), .Y(oclk_1_c));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_3_266_i_m2 (.A(dds_cos[4]), .B(
        sdv_count[1]), .C(dds_sin[4]), .Y(dac1_db_8_3_266_i_m2_net_1));
    CFG4 #( .INIT(16'h1000) )  temp3_49_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_50), .D(N_47), .Y(temp3_49));
    SLE \cnt_freq[3]  (.D(\cnt_freq_s[3] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[3]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  freq3lto8_1 (.A(\data_from_adc[2] [6]), .B(
        \data_from_adc[2] [5]), .C(\data_from_adc[2] [4]), .Y(
        freq3lto8_1_net_1));
    ARI1 #( .INIT(20'h555AA) )  dac_count_1_cry_2 (.A(dac_count[3]), 
        .B(fr_adc_count[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_1_cry_1_net_1), .S(\dac_count_1[3] ), .Y(), .FCO(
        dac_count_1_cry_2_net_1));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_13 (.A(freq_6), .B(
        temp_count[13]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_12_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_13_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[12]  (.A(VCC_net_1), 
        .B(fpga_count[12]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[11]_net_1 ), .S(\fpga_count_s[12] ), .Y(), 
        .FCO(\fpga_count_cry[12]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  GPIO3 (.A(GPIO3_9_net_1), .B(
        GPIO3_8_net_1), .C(GPIO3_7_net_1), .D(GPIO3_6_net_1), .Y(
        GPIO3_c));
    SLE \fpga_count[12]  (.D(\fpga_count_s[12] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[12]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[3]_108 ));
    SLE temp2_csn (.D(\temp_state_i_0[1] ), .CLK(temp_sck_c), .EN(
        temp2_csn_RNO_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_449_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(temp2_csn_c));
    CFG4 #( .INIT(16'h0100) )  freq3lto11 (.A(\data_from_adc[2] [9]), 
        .B(\data_from_adc[2] [11]), .C(\data_from_adc[2] [10]), .D(
        freq3lt11), .Y(freq3));
    SLE \BW_out[11]  (.D(fpga_count[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[11]));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_24 (.A(VCC_net_1), .B(
        temp_count[24]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_23_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_24_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[5]_136 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(N_183), .Y(
        \data_from_adc[2]_96 ));
    SLE \cnt_freq[13]  (.D(\cnt_freq_s[13] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[13]_net_1 ));
    CFG3 #( .INIT(8'h80) )  un1_temp_state28_0_a3_0 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[1]_net_1 ), .C(
        \temp_state[0]_net_1 ), .Y(N_109));
    CFG4 #( .INIT(16'h4000) )  temp2_28_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_48), .Y(temp2_28));
    CFG2 #( .INIT(4'h4) )  \fr_adc_count_5_0_a2[2]  (.A(freq3), .B(
        \un1_data_from_adc[2]_2 ), .Y(\fr_adc_count_5[2] ));
    CFG4 #( .INIT(16'h8000) )  \un1_data_from_adc[2]_1lto11_i_a2_7  (
        .A(\data_from_adc[2] [8]), .B(\data_from_adc[2] [7]), .C(
        \data_from_adc[2] [3]), .D(\data_from_adc[2] [2]), .Y(
        \un1_data_from_adc[2]_1lto11_i_a2_7_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[7]_162 ));
    SLE \temp_count[4]  (.D(\temp_count_s[4] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[4]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIGS2D81[19]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[19]), .D(GND_net_1), .FCI(\temp_count_cry[18] ), .S(
        \temp_count_s[19] ), .Y(), .FCO(\temp_count_cry[19] ));
    SLE \temp_count[10]  (.D(\temp_count_s[10] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[10]));
    SLE \temp3[5]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_39), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[5]));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_29 (.A(VCC_net_1), .B(
        temp_count[29]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_28_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_29_net_1));
    SLE \temp_state[2]  (.D(\temp_state_7[2] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\temp_state[2]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_cry_2 (.A(
        dac_count[2]), .B(fr_adc_count[2]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_fr_adc_count_cry_1_net_1), .S(), .Y(), 
        .FCO(un1_fr_adc_count_cry_2_net_1));
    CFG4 #( .INIT(16'h0040) )  \data_from_adc[6]_0_sqmuxa_3  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ));
    SLE \temp1[3]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_5), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[3]));
    CFG4 #( .INIT(16'h2000) )  temp2_29_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_48), .D(N_47), .Y(temp2_29));
    SLE \fpga_shift_2[2]  (.D(BW_out_c[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[2]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(N_125), .Y(
        \data_from_adc[0]_70 ));
    SLE \data_from_adc[4][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_117 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [0]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_8 (.A(freq_1), .B(
        \cnt_freq[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_7_net_1), .S(), .Y(), .FCO(cnt_freq6_cry_8_net_1)
        );
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIGQGUO1[28]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[28]), .D(GND_net_1), .FCI(\temp_count_cry[27] ), .S(
        \temp_count_s[28] ), .Y(), .FCO(\temp_count_cry[28] ));
    SLE \fpga_shift_2[5]  (.D(BW_out_c[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[5]));
    CFG2 #( .INIT(4'h2) )  \dac_count_3[4]  (.A(\dac_count_1[4] ), .B(
        un1_fr_adc_count_cry_7_net_1), .Y(\dac_count_3[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[7]  (.A(VCC_net_1), .B(
        fpga_count[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[6]_net_1 ), .S(\fpga_count_s[7] ), .Y(), .FCO(
        \fpga_count_cry[7]_net_1 ));
    SLE \temp3[14]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_48), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[14]));
    CFG4 #( .INIT(16'h0C0B) )  temp1_csn_RNO_0 (.A(temp_count_data[4]), 
        .B(\temp_state[0]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(un1_temp_state_8_or));
    CFG4 #( .INIT(16'h6996) )  GPIO5 (.A(GPIO5_14_net_1), .B(
        GPIO5_13_net_1), .C(GPIO5_12_net_1), .D(GPIO5_11_net_1), .Y(
        GPIO5_c));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .Y(\data_from_adc[1]_83 )
        );
    SLE \temp1[11]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_13), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[11]));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_1_cry_5 (.A(
        dac_count[5]), .B(freq_2), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_fr_adc_count_1_cry_4_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_1_cry_5_net_1));
    CFG4 #( .INIT(16'h0400) )  temp3_42_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_50), .Y(temp3_42));
    SLE \temp_count[29]  (.D(\temp_count_s[29] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[29]));
    SLE \data_from_adc[6][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_147 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [6]));
    SLE \temp_count[28]  (.D(\temp_count_s[28] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[28]));
    CFG4 #( .INIT(16'h0100) )  temp1_14_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_49), .Y(temp1_14));
    CFG4 #( .INIT(16'h0C06) )  \cnt_frame_RNO[1]  (.A(
        \cnt_frame[0]_net_1 ), .B(\cnt_frame[1]_net_1 ), .C(N_129), .D(
        N_90), .Y(N_74_i_0));
    SLE \temp2[0]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_18), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[0]));
    SLE \temp2[4]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_22), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[4]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[2]  (.A(
        un13_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[6]_143 ));
    SLE \fpga_count[14]  (.D(\fpga_count_s[14]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[14])
        );
    CFG3 #( .INIT(8'h40) )  \data_from_adc[3]_RNO[0]  (.A(N_82), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(
        \data_from_adc[0]_69_0_0_a2_1 ), .Y(\data_from_adc[3]_105 ));
    SLE \data_from_adc[4][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_122 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [5]));
    ARI1 #( .INIT(20'h45500) )  \cnt_cry_cy[0]  (.A(VCC_net_1), .B(
        un1_cnt_frame_0_sqmuxa_0_net_1), .C(GND_net_1), .D(GND_net_1), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(cnt_cry_cy));
    SLE \fpga_data_receive[5]  (.D(BW_c[5]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[16]  (.A(VCC_net_1), .B(
        \cnt_freq[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[15]_net_1 ), .S(\cnt_freq_s[16] ), .Y(), .FCO(
        \cnt_freq_cry[16]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_27 (.A(VCC_net_1), .B(
        temp_count[27]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_26_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_27_net_1));
    CFG4 #( .INIT(16'h2000) )  temp3_40_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_50), .Y(temp3_40));
    CFG4 #( .INIT(16'h1000) )  temp3_47_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_50), .Y(temp3_47));
    SLE \fr_adc_count[3]  (.D(freq9_i_0_net_1), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fr_adc_count[3]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[25]  (.A(VCC_net_1), .B(
        \cnt_freq[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[24]_net_1 ), .S(\cnt_freq_s[25] ), .Y(), .FCO(
        \cnt_freq_cry[25]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \data_from_adc[2]_RNO[0]  (.A(N_183), .B(
        \data_from_adc[0]_69_0_0_a2_1 ), .C(N_82), .Y(
        \data_from_adc[2]_93 ));
    SLE \data_from_adc[8][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_166 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [1]));
    VCC VCC (.Y(VCC_net_1));
    SLE \temp3[10]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_44), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[10]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[9]  (.A(VCC_net_1), .B(
        fpga_count[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[8]_net_1 ), .S(\fpga_count_s[9] ), .Y(), .FCO(
        \fpga_count_cry[9]_net_1 ));
    CFG2 #( .INIT(4'h1) )  freq3lto3 (.A(\data_from_adc[2] [2]), .B(
        \data_from_adc[2] [3]), .Y(freq3lt8));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(N_185), .C(N_96), .Y(
        \data_from_adc[8]_175 ));
    SLE \data_from_adc[8][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_172 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [7]));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_cry_5 (.A(
        dac_count[5]), .B(freq_2), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_fr_adc_count_cry_4_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_cry_5_net_1));
    CFG4 #( .INIT(16'h0400) )  \data_from_adc[5]_0_sqmuxa_3  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ));
    CFG2 #( .INIT(4'hB) )  un1_cnt_frame_0_sqmuxa_0 (.A(N_130), .B(
        N_90), .Y(un1_cnt_frame_0_sqmuxa_0_net_1));
    SLE \fpga_data_receive[14]  (.D(BW_c[14]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[14]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  \SENSE_DOUT_1_RNO_0[1]  (.A(
        \cnt[5]_net_1 ), .B(\cnt[4]_net_1 ), .C(\cnt[3]_net_1 ), .D(
        N_82), .Y(N_35_i_0));
    SLE \cnt_freq[8]  (.D(\cnt_freq_s[8] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[8]_net_1 ));
    CFG3 #( .INIT(8'h40) )  un20_data_from_adc (.A(\cnt[3]_net_1 ), .B(
        \cnt[1]_net_1 ), .C(GPIO7_c), .Y(un20_data_from_adc_net_1));
    SLE \data_from_adc[3][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_108 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [3]));
    SLE \dac_count[3]  (.D(\dac_count_3[3]_net_1 ), .CLK(BW_clk_c), 
        .EN(clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac_count[3]));
    CFG4 #( .INIT(16'h8000) )  \state_5_i_i_a3_0[0]  (.A(state15), .B(
        SENSE_CS_1_1_sqmuxalt5), .C(\cnt[5]_net_1 ), .D(\cnt[4]_net_1 )
        , .Y(N_130));
    SLE \data_from_adc[4][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_128 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [11]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[1]_88 ));
    SLE \temp1[12]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_14), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[12]));
    CFG4 #( .INIT(16'h6996) )  GPIO5_11 (.A(GPS1_Q1_c), .B(GPS1_Q0_c), 
        .C(GPS1_LD_c), .D(GPS1_I1_c), .Y(GPIO5_11_net_1));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_cry_1 (.A(
        dac_count[1]), .B(fr_adc_count[1]), .C(GND_net_1), .D(
        GND_net_1), .FCI(GND_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_cry_1_net_1));
    SLE \cnt_frame[1]  (.D(N_74_i_0), .CLK(temp_sck_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_frame[1]_net_1 ));
    CFG4 #( .INIT(16'h0200) )  temp2_22_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_48), .Y(temp2_22));
    CFG4 #( .INIT(16'h1000) )  temp2_33_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_48), .D(N_47), .Y(temp2_33));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[7]  (.A(
        un18_data_from_adc_net_1), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[6]_148 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_s[14]  (.A(VCC_net_1), .B(
        fpga_count[14]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[13]_net_1 ), .S(\fpga_count_s[14]_net_1 ), .Y()
        , .FCO());
    SLE \data_from_adc[4][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_121 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [4]));
    SLE \temp3[3]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_37), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[3]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[4]_121 ));
    SLE \data_from_adc[1][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_84 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [3]));
    SLE \cnt_freq[1]  (.D(\cnt_freq_s[1] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  temp2_20_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_48), .Y(temp2_20));
    SLE \BW_out[3]  (.D(fpga_count[3]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[3]));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_1_cry_3 (.A(
        dac_count[3]), .B(fr_adc_count[3]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_fr_adc_count_1_cry_2_net_1), .S(), .Y(), 
        .FCO(un1_fr_adc_count_1_cry_3_net_1));
    CFG4 #( .INIT(16'h4000) )  temp2_27_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_48), .Y(temp2_27));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[27]  (.A(VCC_net_1), .B(
        \cnt_freq[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[26]_net_1 ), .S(\cnt_freq_s[27] ), .Y(), .FCO(
        \cnt_freq_cry[27]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  GPIO3_7 (.A(adc_d0_c[3]), .B(
        adc_d0_c[2]), .C(adc_d0_c[1]), .D(adc_d0_c[0]), .Y(
        GPIO3_7_net_1));
    CFG3 #( .INIT(8'h12) )  \temp_count_data_RNO[1]  (.A(
        temp_count_data[0]), .B(temp_count_data[4]), .C(
        temp_count_data[1]), .Y(N_28_i_0));
    SLE \data_from_adc[2][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_103 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2] [10]));
    ARI1 #( .INIT(20'h42200) )  \cnt_cry[0]  (.A(VCC_net_1), .B(
        GPIO7_c), .C(un1_cnt_frame_0_sqmuxa_0_net_1), .D(GND_net_1), 
        .FCI(cnt_cry_cy), .S(\cnt_s[0] ), .Y(), .FCO(
        \cnt_cry[0]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[3]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(\data_from_adc[3]_0_sqmuxa_3_net_1 ), 
        .Y(\data_from_adc[3]_111 ));
    SLE \data_from_adc[4][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_126 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [9]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[7]  (.A(VCC_net_1), .B(
        \cnt_freq[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[6]_net_1 ), .S(\cnt_freq_s[7] ), .Y(), .FCO(
        \cnt_freq_cry[7]_net_1 ));
    SLE \temp_count_data[4]  (.D(N_7_i_0), .CLK(temp_sck_c), .EN(
        un1_temp_state28_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count_data[4]));
    SLE \dac1_db[6]  (.D(dac1_db_8_0_296_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[6]));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[2]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(N_183), .Y(\data_from_adc[2]_99 ));
    SLE \temp1[1]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_3), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[1]));
    SLE clk_dac1 (.D(clk_dac1_2_net_1), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dac1_clk_c));
    SLE \cnt_freq[7]  (.D(\cnt_freq_s[7] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[7]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI771EJ1[25]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[25]), .D(GND_net_1), .FCI(\temp_count_cry[24] ), .S(
        \temp_count_s[25] ), .Y(), .FCO(\temp_count_cry[25] ));
    SLE \temp_count[7]  (.D(\temp_count_s[7] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[7]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(N_185), .C(N_96), .Y(
        \data_from_adc[8]_169 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIIP6KS1[30]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[30]), .D(GND_net_1), .FCI(\temp_count_cry[29] ), .S(
        \temp_count_s[30] ), .Y(), .FCO(\temp_count_cry[30] ));
    CFG4 #( .INIT(16'h2000) )  temp1_7_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_49), .Y(temp1_7));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[4]  (.A(VCC_net_1), .B(
        \cnt_freq[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[3]_net_1 ), .S(\cnt_freq_s[4] ), .Y(), .FCO(
        \cnt_freq_cry[4]_net_1 ));
    SLE \freq[18]  (.D(\un1_data_from_adc[2]_2 ), .CLK(temp_sck_c), 
        .EN(\un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_11));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[4]_126 ));
    CFG4 #( .INIT(16'h00AE) )  \cnt_frame_0_0[3]  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame_0_0_a3_0_1_0[3]_net_1 ), 
        .C(N_105), .D(N_129), .Y(\cnt_frame_0_0[3]_net_1 ));
    CFG2 #( .INIT(4'h7) )  temp_count_data_n3_i_o2 (.A(
        temp_count_data[0]), .B(temp_count_data[1]), .Y(N_73));
    CFG4 #( .INIT(16'h0200) )  temp3_38_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_50), .Y(temp3_38));
    SLE \data_from_adc[1][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_92 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [11]));
    SLE \temp_count[5]  (.D(\temp_count_s[5] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[5]));
    SLE \temp_count[0]  (.D(\temp_count_s[0] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[0]));
    SLE \temp_count[31]  (.D(\temp_count_s[31] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[31]));
    SLE \data_from_adc[4][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_125 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [8]));
    SLE \temp3[2]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_36), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[2]));
    CFG4 #( .INIT(16'h4414) )  \temp_count_data_RNO[3]  (.A(
        temp_count_data[4]), .B(temp_count_data[3]), .C(
        temp_count_data[2]), .D(N_73), .Y(N_9_i_0));
    SLE \fpga_data_receive[3]  (.D(BW_c[3]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[3]_net_1 ));
    SLE \dac1_db[7]  (.D(dac1_db_8_1_286_i_m2_net_1), .CLK(BW_clk_c), 
        .EN(\sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        dac1_db_c[7]));
    SLE \temp2[6]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_24), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[6]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[29]  (.A(VCC_net_1), .B(
        \cnt_freq[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[28]_net_1 ), .S(\cnt_freq_s[29] ), .Y(), .FCO(
        \cnt_freq_cry[29]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[7]_154 ));
    SLE \data_from_adc[3][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_111 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [6]));
    SLE \data_from_adc[6][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_142 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [1]));
    ARI1 #( .INIT(20'h44400) )  \cnt_s[5]  (.A(VCC_net_1), .B(
        un1_cnt_frame_0_sqmuxa_0_net_1), .C(\cnt[5]_net_1 ), .D(
        GND_net_1), .FCI(\cnt_cry[4]_net_1 ), .S(\cnt_s[5]_net_1 ), .Y(
        ), .FCO());
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_39 (.A(
        \fpga_data_receive[3]_net_1 ), .B(fpga_shift_2[2]), .C(
        fpga_shift_2[3]), .D(\fpga_data_receive[2]_net_1 ), .FCI(
        \fpga_flag4_0_data_tmp[0] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[1] ));
    CFG4 #( .INIT(16'h2000) )  temp3_39_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_50), .Y(temp3_39));
    SLE \temp_count[19]  (.D(\temp_count_s[19] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[19]));
    SLE \fpga_data_receive[12]  (.D(BW_c[12]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[12]_net_1 ));
    SLE \temp_count[18]  (.D(\temp_count_s[18] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[18]));
    CFG4 #( .INIT(16'h4000) )  temp1_9_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_49), .D(N_47), .Y(temp1_9));
    SLE \fpga_count[11]  (.D(\fpga_count_s[11] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[11]));
    SLE \data_from_adc[6][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_148 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [7]));
    SLE \data_from_adc[0][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_69 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [0]));
    SLE clk_dac2_inst_1 (.D(sdv_count[0]), .CLK(BW_clk_c), .EN(
        sdv_count[1]), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(clk_dac2));
    CFG4 #( .INIT(16'h1000) )  temp2_31_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_48), .Y(temp2_31));
    CFG4 #( .INIT(16'h4000) )  temp3_44_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_50), .Y(temp3_44));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_0_296_i_m2 (.A(dds_cos[1]), .B(
        sdv_count[1]), .C(dds_sin[1]), .Y(dac1_db_8_0_296_i_m2_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[5]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[5]_132 ));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_cry_3 (.A(
        dac_count[3]), .B(fr_adc_count[3]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_fr_adc_count_cry_2_net_1), .S(), .Y(), 
        .FCO(un1_fr_adc_count_cry_3_net_1));
    SLE \data_from_adc[1][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_87 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [6]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[8]_RNO[9]  (.A(
        un20_data_from_adc_net_1), .B(N_185), .C(N_96), .Y(
        \data_from_adc[8]_174 ));
    SLE \data_from_adc[0][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_74 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [5]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[5]  (.A(_decfrac4), 
        .B(N_96), .C(N_125), .Y(\data_from_adc[0]_74 ));
    SLE \cnt[1]  (.D(\cnt_s[1] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[1]_net_1 ));
    CFG4 #( .INIT(16'hC8CC) )  \un1_data_from_adc[2]_2lto11_i  (.A(
        \data_from_adc[2] [9]), .B(\data_from_adc[2] [11]), .C(
        \data_from_adc[2] [10]), .D(\un1_data_from_adc[2]_2lt10 ), .Y(
        \un1_data_from_adc[2]_2_i_0 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9QGHR[12]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[12]), .D(GND_net_1), .FCI(\temp_count_cry[11] ), .S(
        \temp_count_s[12] ), .Y(), .FCO(\temp_count_cry[12] ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[6]  (.A(VCC_net_1), .B(
        fpga_count[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[5]_net_1 ), .S(\fpga_count_s[6] ), .Y(), .FCO(
        \fpga_count_cry[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[13]  (.A(VCC_net_1), .B(
        \cnt_freq[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[12]_net_1 ), .S(\cnt_freq_s[13] ), .Y(), .FCO(
        \cnt_freq_cry[13]_net_1 ));
    SLE \data_from_adc[8][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[8]_167 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[8] [2]));
    SLE \BW_out[12]  (.D(fpga_count[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[12]));
    CFG4 #( .INIT(16'h0002) )  \data_from_adc[8]_0_sqmuxa_0_a2  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[1]_net_1 ), .D(\cnt_frame[0]_net_1 ), .Y(N_185));
    SLE \temp2[15]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_33), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[15]));
    SLE GPIO16 (.D(N_13_i_0), .CLK(temp_sck_c), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(GPIO16_c));
    CFG4 #( .INIT(16'h2000) )  temp2_24_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_48), .Y(temp2_24));
    SLE \fpga_count[7]  (.D(\fpga_count_s[7] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[7]));
    SLE \temp_count[24]  (.D(\temp_count_s[24] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[24]));
    CFG4 #( .INIT(16'h8B33) )  \temp_state_7_2_0_.m7_am  (.A(GPIO11_c), 
        .B(\temp_state[1]_net_1 ), .C(temp_count_data[4]), .D(
        \temp_state[0]_net_1 ), .Y(m7_am));
    ARI1 #( .INIT(20'h555AA) )  dac_count_1_cry_4 (.A(dac_count[5]), 
        .B(freq_2), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_1_cry_3_net_1), .S(\dac_count_1[5] ), .Y(), .FCO(
        dac_count_1_cry_4_net_1));
    SLE \cnt_freq[29]  (.D(\cnt_freq_s[29] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[29]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[10]  (.A(
        un21_data_from_adc_net_1), .B(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[7]_163 ));
    SLE \cnt_frame[0]  (.D(N_76_i_0), .CLK(temp_sck_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_frame[0]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[5]_RNO[0]  (.A(N_82), .B(
        \data_from_adc[5]_0_sqmuxa_3_net_1 ), .C(
        \data_from_adc[0]_69_0_0_a2_1 ), .Y(\data_from_adc[5]_129 ));
    SLE \data_from_adc[0][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_73 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [4]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[4]  (.A(VCC_net_1), .B(
        fpga_count[4]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[3]_net_1 ), .S(\fpga_count_s[4] ), .Y(), .FCO(
        \fpga_count_cry[4]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  temp2_18_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_48), .Y(temp2_18));
    CFG2 #( .INIT(4'hE) )  temp1_csn_RNO (.A(temp_state26), .B(
        un1_temp_state_8_or), .Y(temp1_csn_RNO_net_1));
    SLE \data_from_adc[5][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_129 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [0]));
    SLE \fpga_shift_2[9]  (.D(BW_out_c[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[9]));
    CFG4 #( .INIT(16'h8000) )  temp3_37_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_50), .D(N_47), .Y(temp3_37));
    SLE \temp_count_data[1]  (.D(N_28_i_0), .CLK(temp_sck_c), .EN(
        un1_temp_state28_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count_data[1]));
    SLE \BW_out[7]  (.D(fpga_count[7]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[7]));
    SLE \BW_out[4]  (.D(fpga_count[4]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[4]));
    SLE \temp3[4]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_38), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[4]));
    SLE \cnt[2]  (.D(\cnt_s[2] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[2]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNILDBPQ1[29]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[29]), .D(GND_net_1), .FCI(\temp_count_cry[28] ), .S(
        \temp_count_s[29] ), .Y(), .FCO(\temp_count_cry[29] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[1]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .Y(\data_from_adc[1]_84 )
        );
    CFG4 #( .INIT(16'h8000) )  temp2_19_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_48), .Y(temp2_19));
    SLE \data_from_adc[0][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_78 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [9]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[6]  (.A(VCC_net_1), .B(
        \cnt_freq[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[5]_net_1 ), .S(\cnt_freq_s[6] ), .Y(), .FCO(
        \cnt_freq_cry[6]_net_1 ));
    SLE \cnt_freq[4]  (.D(\cnt_freq_s[4] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[4]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[3]  (.A(
        un14_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[6]_144 ));
    SLE \data_from_adc[5][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_134 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [5]));
    CFG3 #( .INIT(8'h08) )  \data_from_adc[0]_RNO[8]  (.A(N_125), .B(
        N_168), .C(N_82), .Y(\data_from_adc[0]_77 ));
    CFG4 #( .INIT(16'h8000) )  temp1_4_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_49), .Y(temp1_4));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_25 (.A(VCC_net_1), .B(
        \cnt_freq[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_24_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_25_net_1));
    SLE \cnt_freq[19]  (.D(\cnt_freq_s[19] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[19]_net_1 ));
    CFG4 #( .INIT(16'h000E) )  \SENSE_DOUT_1_RNO[1]  (.A(N_714), .B(
        N_105), .C(\SENSE_DOUT_2_1_u_i_0[1]_net_1 ), .D(
        \SENSE_DOUT_2_1_u_i_1[1]_net_1 ), .Y(N_37_i_0));
    CFG4 #( .INIT(16'hCECC) )  \SENSE_DOUT_2_1_u_i_1[1]  (.A(N_170), 
        .B(N_125), .C(GPIO7_c), .D(
        \SENSE_DOUT_2_1_u_i_a3_3_0[1]_net_1 ), .Y(
        \SENSE_DOUT_2_1_u_i_1[1]_net_1 ));
    SLE \fpga_data_receive[10]  (.D(BW_c[10]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[10]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_1_cry_1 (.A(
        dac_count[1]), .B(fr_adc_count[1]), .C(GND_net_1), .D(
        GND_net_1), .FCI(GND_net_1), .S(), .Y(), .FCO(
        un1_fr_adc_count_1_cry_1_net_1));
    CFG4 #( .INIT(16'h002E) )  \state_RNO[1]  (.A(\state[1]_net_1 ), 
        .B(\state[0]_net_1 ), .C(\cnt_frame[3]_net_1 ), .D(N_130), .Y(
        N_40_i_0));
    CFG3 #( .INIT(8'h40) )  temp_state26_0_a3 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[1]_net_1 ), .C(
        \temp_state[0]_net_1 ), .Y(temp_state26));
    SLE \data_from_adc[3][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_106 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [1]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[3]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(
        \data_from_adc[3]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[3]_109 ));
    CFG4 #( .INIT(16'h6996) )  GPIO5_13 (.A(adc_of_c), .B(adc_oen_c), 
        .C(adc_clk_c), .D(GPS_I1_c), .Y(GPIO5_13_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[0]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(N_125), .C(N_96), .Y(
        \data_from_adc[0]_80 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_16 (.A(freq_1), .B(
        temp_count[16]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_15_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_16_net_1));
    ARI1 #( .INIT(20'h555AA) )  un1_fr_adc_count_1_cry_4 (.A(
        dac_count[4]), .B(fr_adc_count[2]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_fr_adc_count_1_cry_3_net_1), .S(), .Y(), 
        .FCO(un1_fr_adc_count_1_cry_4_net_1));
    CFG4 #( .INIT(16'h1000) )  temp1_15_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_52), .D(N_49), .Y(temp1_15));
    SLE \data_from_adc[3][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[3]_112 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[3] [7]));
    SLE \data_from_adc[7][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_164 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [11]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[4]_RNO[1]  (.A(
        un12_data_from_adc_net_1), .B(N_96), .C(
        \data_from_adc[4]_0_sqmuxa_3_net_1 ), .Y(
        \data_from_adc[4]_118 ));
    CFG4 #( .INIT(16'h1000) )  temp1_16_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_49), .Y(temp1_16));
    CFG3 #( .INIT(8'h04) )  un22_data_from_adc (.A(\cnt[3]_net_1 ), .B(
        \cnt[2]_net_1 ), .C(\cnt[1]_net_1 ), .Y(
        un22_data_from_adc_net_1));
    SLE \fpga_count[10]  (.D(\fpga_count_s[10] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[10]));
    CFG4 #( .INIT(16'h4000) )  \data_from_adc[5]_RNO[6]  (.A(GPIO7_c), 
        .B(N_170), .C(N_168), .D(\data_from_adc[5]_0_sqmuxa_3_net_1 ), 
        .Y(\data_from_adc[5]_135 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[4]  (.A(
        un15_data_from_adc_net_1), .B(N_183), .C(N_96), .Y(
        \data_from_adc[2]_97 ));
    CFG4 #( .INIT(16'h1000) )  temp2_32_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_51), .D(N_48), .Y(temp2_32));
    SLE \fpga_shift_2[6]  (.D(BW_out_c[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[6]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_30 (.A(VCC_net_1), .B(
        \cnt_freq[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_29_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_30_net_1));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_18 (.A(freq_11), .B(
        temp_count[18]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_17_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_18_net_1));
    SLE \cnt_freq[6]  (.D(\cnt_freq_s[6] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[6]_net_1 ));
    SLE \data_from_adc[7][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_153 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [0]));
    SLE \data_from_adc[0][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_77 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [8]));
    SLE \fpga_count[2]  (.D(\fpga_count_s[2] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_count[2]));
    SLE \data_from_adc[5][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_133 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [4]));
    SLE \data_from_adc[0][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[0]_79 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[0] [10]));
    CFG2 #( .INIT(4'h6) )  GPIO3_6 (.A(adc_d0_c[12]), .B(adc_d0_c[13]), 
        .Y(GPIO3_6_net_1));
    SLE \data_from_adc[6][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[6]_143 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[6] [2]));
    SLE \data_from_adc[4][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[4]_120 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[4] [3]));
    SLE \data_from_adc[1][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_82 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [1]));
    ARI1 #( .INIT(20'h4AA00) )  fpga_count_s_530 (.A(VCC_net_1), .B(
        fpga_count[0]), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(fpga_count_s_530_FCO));
    CFG1 #( .INIT(2'h1) )  \sdv_count_RNI847F[0]  (.A(sdv_count[0]), 
        .Y(\sdv_count_i_0[0] ));
    SLE GPIO14 (.D(fpga_flag_net_1), .CLK(BW_clk_c_i_0), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(GPIO14_c));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[1]_RNO[0]  (.A(N_82), .B(
        \data_from_adc[1]_0_sqmuxa_3_net_1 ), .C(
        \data_from_adc[0]_69_0_0_a2_1 ), .Y(\data_from_adc[1]_81 ));
    CFG3 #( .INIT(8'hD8) )  \temp_state_7_2_0_.m7_ns  (.A(
        \temp_state[2]_net_1 ), .B(m7_bm), .C(m7_am), .Y(
        \temp_state_7[0] ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[5]  (.A(VCC_net_1), .B(
        \cnt_freq[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[4]_net_1 ), .S(\cnt_freq_s[5] ), .Y(), .FCO(
        \cnt_freq_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  temp2_30_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_73), .D(N_48), .Y(temp2_30));
    SLE \data_from_adc[1][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[1]_88 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[1] [7]));
    SLE \temp_count_data[2]  (.D(N_11_i_0), .CLK(temp_sck_c), .EN(
        un1_temp_state28_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count_data[2]));
    SLE \fpga_shift_2[14]  (.D(BW_out_c[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(fpga_shift_2[14]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI2MNTJ[8]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[8]), .D(
        GND_net_1), .FCI(\temp_count_cry[7] ), .S(\temp_count_s[8] ), 
        .Y(), .FCO(\temp_count_cry[8] ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[3]  (.A(VCC_net_1), .B(
        fpga_count[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[2]_net_1 ), .S(\fpga_count_s[3] ), .Y(), .FCO(
        \fpga_count_cry[3]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  dac1_db_8_5_246_i_m2 (.A(dds_cos[6]), .B(
        sdv_count[1]), .C(dds_sin[6]), .Y(dac1_db_8_5_246_i_m2_net_1));
    CFG3 #( .INIT(8'h40) )  \data_from_adc[6]_RNO[0]  (.A(N_82), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(
        \data_from_adc[0]_69_0_0_a2_1 ), .Y(\data_from_adc[6]_141 ));
    CFG4 #( .INIT(16'hC080) )  \data_from_adc[2]_0_sqmuxa_0_a2_3_RNO  
        (.A(GPIO7_c), .B(data_m1_e_0_1), .C(\cnt[2]_net_1 ), .D(
        \cnt[1]_net_1 ), .Y(
        \data_from_adc[2]_0_sqmuxa_0_a2_3_RNO_net_1 ));
    SLE \data_from_adc[7][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[7]_158 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[7] [5]));
    SLE \freq[8]  (.D(freq3), .CLK(temp_sck_c), .EN(
        \un1_data_from_adc[2]_1_i_i_0 ), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(freq_1));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_15 (.A(freq_0), .B(
        \cnt_freq[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_14_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_15_net_1));
    SLE \data_from_adc[5][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_138 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [9]));
    SLE \data_from_adc[5][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[5]_139 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[5] [10]));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_25 (.A(VCC_net_1), .B(
        temp_count[25]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_24_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_25_net_1));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_21 (.A(
        \fpga_data_receive[9]_net_1 ), .B(fpga_shift_2[8]), .C(
        fpga_shift_2[9]), .D(\fpga_data_receive[8]_net_1 ), .FCI(
        \fpga_flag4_0_data_tmp[3] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[4] ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[6]_RNO[11]  (.A(
        un22_data_from_adc_net_1), .B(
        \data_from_adc[6]_0_sqmuxa_3_net_1 ), .C(N_96), .Y(
        \data_from_adc[6]_152 ));
    SLE \cnt_freq[21]  (.D(\cnt_freq_s[21] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[21]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[7]_RNO[5]  (.A(
        \data_from_adc[7]_0_sqmuxa_3_net_1 ), .B(_decfrac4), .C(N_96), 
        .Y(\data_from_adc[7]_158 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[10]  (.A(VCC_net_1), 
        .B(fpga_count[10]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[9]_net_1 ), .S(\fpga_count_s[10] ), .Y(), .FCO(
        \fpga_count_cry[10]_net_1 ));
    
endmodule


module b5_nvmFL_1131s_x(
       b4_nUAi,
       IICE_comm2iice,
       b4_PLyF,
       b7_PSyi3wy,
       b8_PSyiBgYG
    );
output [1129:0] b4_nUAi;
input  [11:10] IICE_comm2iice;
input  b4_PLyF;
output b7_PSyi3wy;
input  b8_PSyiBgYG;

    wire VCC_net_1, b6_OKctIF4_net_1, GND_net_1;
    
    SLE \b6_OKctIF[789]  (.D(b4_nUAi[340]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[341]));
    SLE \b6_OKctIF[310]  (.D(b4_nUAi[819]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[820]));
    SLE \b6_OKctIF[247]  (.D(b4_nUAi[882]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[883]));
    SLE \b6_OKctIF[393]  (.D(b4_nUAi[736]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[737]));
    SLE \b6_OKctIF[876]  (.D(b4_nUAi[253]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[254]));
    SLE \b6_OKctIF[1047]  (.D(b4_nUAi[82]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[83]));
    SLE \b6_OKctIF[297]  (.D(b4_nUAi[832]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[833]));
    SLE \b6_OKctIF[235]  (.D(b4_nUAi[894]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[895]));
    SLE \b6_OKctIF[465]  (.D(b4_nUAi[664]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[665]));
    SLE \b6_OKctIF[430]  (.D(b4_nUAi[699]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[700]));
    SLE \b6_OKctIF[332]  (.D(b4_nUAi[797]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[798]));
    SLE \b6_OKctIF[862]  (.D(b4_nUAi[267]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[268]));
    SLE \b6_OKctIF[75]  (.D(b4_nUAi[1054]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1055]));
    SLE \b6_OKctIF[1043]  (.D(b4_nUAi[86]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[87]));
    SLE \b6_OKctIF[216]  (.D(b4_nUAi[913]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[914]));
    SLE \b6_OKctIF[70]  (.D(b4_nUAi[1059]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1060]));
    SLE \b6_OKctIF[1019]  (.D(b4_nUAi[110]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[111]));
    SLE \b6_OKctIF[1123]  (.D(b4_nUAi[6]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[7]));
    SLE \b6_OKctIF[666]  (.D(b4_nUAi[463]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[464]));
    SLE \b6_OKctIF[205]  (.D(b4_nUAi[924]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[925]));
    SLE \b6_OKctIF[471]  (.D(b4_nUAi[658]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[659]));
    SLE \b6_OKctIF[400]  (.D(b4_nUAi[729]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[730]));
    SLE \b6_OKctIF[414]  (.D(b4_nUAi[715]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[716]));
    SLE \b6_OKctIF[883]  (.D(b4_nUAi[246]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[247]));
    SLE \b6_OKctIF[766]  (.D(b4_nUAi[363]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[364]));
    SLE \b6_OKctIF[552]  (.D(b4_nUAi[577]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[578]));
    SLE \b6_OKctIF[467]  (.D(b4_nUAi[662]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[663]));
    SLE \b6_OKctIF[328]  (.D(b4_nUAi[801]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[802]));
    SLE \b6_OKctIF[302]  (.D(b4_nUAi[827]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[828]));
    SLE \b6_OKctIF[27]  (.D(b4_nUAi[1102]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1103]));
    SLE \b6_OKctIF[628]  (.D(b4_nUAi[501]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[502]));
    SLE \b6_OKctIF[542]  (.D(b4_nUAi[587]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[588]));
    SLE \b6_OKctIF[685]  (.D(b4_nUAi[444]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[445]));
    SLE \b6_OKctIF[365]  (.D(b4_nUAi[764]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[765]));
    SLE \b6_OKctIF[177]  (.D(b4_nUAi[952]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[953]));
    SLE \b6_OKctIF[921]  (.D(b4_nUAi[208]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[209]));
    SLE \b6_OKctIF[58]  (.D(b4_nUAi[1071]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1072]));
    SLE \b6_OKctIF[24]  (.D(b4_nUAi[1105]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1106]));
    SLE \b6_OKctIF[1024]  (.D(b4_nUAi[105]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[106]));
    SLE \b6_OKctIF[592]  (.D(b4_nUAi[537]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[538]));
    SLE \b6_OKctIF[180]  (.D(b4_nUAi[949]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[950]));
    SLE \b6_OKctIF[111]  (.D(b4_nUAi[1018]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1019]));
    SLE \b6_OKctIF[651]  (.D(b4_nUAi[478]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[479]));
    SLE \b6_OKctIF[158]  (.D(b4_nUAi[971]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[972]));
    SLE \b6_OKctIF[1122]  (.D(b4_nUAi[7]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[8]));
    SLE \b6_OKctIF[29]  (.D(b4_nUAi[1100]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1101]));
    SLE \b6_OKctIF[857]  (.D(b4_nUAi[272]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[273]));
    SLE \b6_OKctIF[641]  (.D(b4_nUAi[488]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[489]));
    SLE \b6_OKctIF[623]  (.D(b4_nUAi[506]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[507]));
    SLE \b6_OKctIF[319]  (.D(b4_nUAi[810]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[811]));
    SLE \b6_OKctIF[262]  (.D(b4_nUAi[867]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[868]));
    SLE \b6_OKctIF[148]  (.D(b4_nUAi[981]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[982]));
    SLE \b6_OKctIF[165]  (.D(b4_nUAi[964]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[965]));
    SLE \b6_OKctIF[847]  (.D(b4_nUAi[282]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[283]));
    SLE \b6_OKctIF[123]  (.D(b4_nUAi[1006]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1007]));
    SLE \b6_OKctIF[566]  (.D(b4_nUAi[563]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[564]));
    SLE \b6_OKctIF[456]  (.D(b4_nUAi[673]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[674]));
    SLE \b6_OKctIF[734]  (.D(b4_nUAi[395]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[396]));
    SLE \b6_OKctIF[691]  (.D(b4_nUAi[438]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[439]));
    SLE \b6_OKctIF[198]  (.D(b4_nUAi[931]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[932]));
    SLE \b6_OKctIF[725]  (.D(b4_nUAi[404]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[405]));
    SLE \b6_OKctIF[51]  (.D(b4_nUAi[1078]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1079]));
    SLE \b6_OKctIF[446]  (.D(b4_nUAi[683]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[684]));
    SLE \b6_OKctIF[897]  (.D(b4_nUAi[232]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[233]));
    SLE \b6_OKctIF[77]  (.D(b4_nUAi[1052]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1053]));
    SLE \b6_OKctIF[136]  (.D(b4_nUAi[993]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[994]));
    SLE \b6_OKctIF[580]  (.D(b4_nUAi[549]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[550]));
    SLE \b6_OKctIF[704]  (.D(b4_nUAi[425]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[426]));
    SLE \b6_OKctIF[288]  (.D(b4_nUAi[841]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[842]));
    SLE \b6_OKctIF[757]  (.D(b4_nUAi[372]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[373]));
    SLE \b6_OKctIF[74]  (.D(b4_nUAi[1055]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1056]));
    SLE \b6_OKctIF[496]  (.D(b4_nUAi[633]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[634]));
    SLE \b6_OKctIF[1040]  (.D(b4_nUAi[89]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[90]));
    SLE \b6_OKctIF[815]  (.D(b4_nUAi[314]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[315]));
    SLE \b6_OKctIF[829]  (.D(b4_nUAi[300]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[301]));
    SLE \b6_OKctIF[747]  (.D(b4_nUAi[382]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[383]));
    SLE \b6_OKctIF[106]  (.D(b4_nUAi[1023]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1024]));
    SLE \b6_OKctIF[733]  (.D(b4_nUAi[396]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[397]));
    SLE \b6_OKctIF[915]  (.D(b4_nUAi[214]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[215]));
    SLE \b6_OKctIF[929]  (.D(b4_nUAi[200]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[201]));
    SLE \b6_OKctIF[1065]  (.D(b4_nUAi[64]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[65]));
    SLE \b6_OKctIF[567]  (.D(b4_nUAi[562]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[563]));
    SLE \b6_OKctIF[838]  (.D(b4_nUAi[291]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[292]));
    SLE \b6_OKctIF[79]  (.D(b4_nUAi[1050]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1051]));
    SLE \b6_OKctIF[164]  (.D(b4_nUAi[965]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[966]));
    SLE \b6_OKctIF[558]  (.D(b4_nUAi[571]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[572]));
    SLE \b6_OKctIF[233]  (.D(b4_nUAi[896]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[897]));
    SLE \b6_OKctIF[48]  (.D(b4_nUAi[1081]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1082]));
    SLE \b6_OKctIF[797]  (.D(b4_nUAi[332]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[333]));
    SLE \b6_OKctIF[703]  (.D(b4_nUAi[426]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[427]));
    SLE \b6_OKctIF[548]  (.D(b4_nUAi[581]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[582]));
    SLE \b6_OKctIF[927]  (.D(b4_nUAi[202]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[203]));
    SLE \b6_OKctIF[351]  (.D(b4_nUAi[778]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[779]));
    SLE \b6_OKctIF[808]  (.D(b4_nUAi[321]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[322]));
    SLE \b6_OKctIF[357]  (.D(b4_nUAi[772]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[773]));
    SLE \b6_OKctIF[583]  (.D(b4_nUAi[546]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[547]));
    SLE \b6_OKctIF[203]  (.D(b4_nUAi[926]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[927]));
    SLE \b6_OKctIF[824]  (.D(b4_nUAi[305]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[306]));
    SLE \b6_OKctIF[535]  (.D(b4_nUAi[594]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[595]));
    SLE \b6_OKctIF[341]  (.D(b4_nUAi[788]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[789]));
    SLE \b6_OKctIF[482]  (.D(b4_nUAi[647]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[648]));
    SLE \b6_OKctIF[598]  (.D(b4_nUAi[531]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[532]));
    SLE \b6_OKctIF[347]  (.D(b4_nUAi[782]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[783]));
    SLE \b6_OKctIF[680]  (.D(b4_nUAi[449]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[450]));
    SLE \b6_OKctIF[428]  (.D(b4_nUAi[701]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[702]));
    SLE \b6_OKctIF[483]  (.D(b4_nUAi[646]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[647]));
    SLE \b6_OKctIF[215]  (.D(b4_nUAi[914]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[915]));
    SLE \b6_OKctIF[410]  (.D(b4_nUAi[719]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[720]));
    SLE \b6_OKctIF[571]  (.D(b4_nUAi[558]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[559]));
    SLE \b6_OKctIF[312]  (.D(b4_nUAi[817]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[818]));
    SLE \b6_OKctIF[505]  (.D(b4_nUAi[624]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[625]));
    SLE \b6_OKctIF[391]  (.D(b4_nUAi[738]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[739]));
    SLE \b6_OKctIF[627]  (.D(b4_nUAi[502]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[503]));
    SLE \b6_OKctIF[397]  (.D(b4_nUAi[732]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[733]));
    SLE \b6_OKctIF[41]  (.D(b4_nUAi[1088]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1089]));
    SLE \b6_OKctIF[230]  (.D(b4_nUAi[899]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[900]));
    SLE \b6_OKctIF[936]  (.D(b4_nUAi[193]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[194]));
    SLE \b6_OKctIF[953]  (.D(b4_nUAi[176]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[177]));
    SLE \b6_OKctIF[289]  (.D(b4_nUAi[840]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[841]));
    SLE \b6_OKctIF[354]  (.D(b4_nUAi[775]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[776]));
    SLE \b6_OKctIF[1021]  (.D(b4_nUAi[108]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[109]));
    SLE \b6_OKctIF[479]  (.D(b4_nUAi[650]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[651]));
    SLE \b6_OKctIF[943]  (.D(b4_nUAi[186]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[187]));
    SLE \b6_OKctIF[376]  (.D(b4_nUAi[753]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[754]));
    SLE \b6_OKctIF[368]  (.D(b4_nUAi[761]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[762]));
    SLE \b6_OKctIF[344]  (.D(b4_nUAi[785]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[786]));
    SLE \b6_OKctIF[200]  (.D(b4_nUAi[929]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[930]));
    SLE \b6_OKctIF[1088]  (.D(b4_nUAi[41]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[42]));
    SLE \b6_OKctIF[906]  (.D(b4_nUAi[223]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[224]));
    SLE \b6_OKctIF[668]  (.D(b4_nUAi[461]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[462]));
    SLE \b6_OKctIF[836]  (.D(b4_nUAi[293]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[294]));
    SLE \b6_OKctIF[993]  (.D(b4_nUAi[136]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[137]));
    SLE \b6_OKctIF[961]  (.D(b4_nUAi[168]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[169]));
    SLE \b6_OKctIF[394]  (.D(b4_nUAi[735]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[736]));
    SLE \b6_OKctIF[56]  (.D(b4_nUAi[1073]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1074]));
    SLE \b6_OKctIF[806]  (.D(b4_nUAi[323]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[324]));
    SLE \b6_OKctIF[759]  (.D(b4_nUAi[370]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[371]));
    SLE \b6_OKctIF[431]  (.D(b4_nUAi[698]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[699]));
    SLE \b6_OKctIF[1029]  (.D(b4_nUAi[100]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[101]));
    SLE \b6_OKctIF[749]  (.D(b4_nUAi[380]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[381]));
    SLE \b6_OKctIF[974]  (.D(b4_nUAi[155]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[156]));
    SLE \b6_OKctIF[728]  (.D(b4_nUAi[401]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[402]));
    SLE \b6_OKctIF[663]  (.D(b4_nUAi[466]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[467]));
    SLE \b6_OKctIF[182]  (.D(b4_nUAi[947]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[948]));
    SLE \b6_OKctIF[782]  (.D(b4_nUAi[347]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[348]));
    SLE \b6_OKctIF[714]  (.D(b4_nUAi[415]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[416]));
    SLE \b6_OKctIF[401]  (.D(b4_nUAi[728]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[729]));
    SLE \b6_OKctIF[163]  (.D(b4_nUAi[966]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[967]));
    SLE \b6_OKctIF[137]  (.D(b4_nUAi[992]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[993]));
    SLE \b6_OKctIF[629]  (.D(b4_nUAi[500]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[501]));
    SLE \b6_OKctIF[1094]  (.D(b4_nUAi[35]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[36]));
    SLE \b6_OKctIF[870]  (.D(b4_nUAi[259]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[260]));
    SLE \b6_OKctIF[799]  (.D(b4_nUAi[330]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[331]));
    SLE \b6_OKctIF[1032]  (.D(b4_nUAi[97]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[98]));
    SLE \b6_OKctIF[116]  (.D(b4_nUAi[1013]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1014]));
    SLE \b6_OKctIF[765]  (.D(b4_nUAi[364]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[365]));
    SLE \b6_OKctIF[920]  (.D(b4_nUAi[209]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[210]));
    SLE \b6_OKctIF[853]  (.D(b4_nUAi[276]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[277]));
    SLE \b6_OKctIF[107]  (.D(b4_nUAi[1022]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1023]));
    SLE \b6_OKctIF[1036]  (.D(b4_nUAi[93]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[94]));
    SLE \b6_OKctIF[843]  (.D(b4_nUAi[286]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[287]));
    SLE \b6_OKctIF[713]  (.D(b4_nUAi[416]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[417]));
    SLE \b6_OKctIF[655]  (.D(b4_nUAi[474]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[475]));
    SLE \b6_OKctIF[869]  (.D(b4_nUAi[260]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[261]));
    SLE \b6_OKctIF[821]  (.D(b4_nUAi[308]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[309]));
    SLE \b6_OKctIF[485]  (.D(b4_nUAi[644]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[645]));
    SLE \b6_OKctIF[882]  (.D(b4_nUAi[247]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[248]));
    SLE \b6_OKctIF[818]  (.D(b4_nUAi[311]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[312]));
    SLE \b6_OKctIF[213]  (.D(b4_nUAi[916]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[917]));
    SLE \b6_OKctIF[969]  (.D(b4_nUAi[160]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[161]));
    SLE \b6_OKctIF[645]  (.D(b4_nUAi[484]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[485]));
    SLE \b6_OKctIF[1072]  (.D(b4_nUAi[57]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[58]));
    SLE \b6_OKctIF[893]  (.D(b4_nUAi[236]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[237]));
    SLE \b6_OKctIF[150]  (.D(b4_nUAi[979]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[980]));
    GND GND (.Y(GND_net_1));
    SLE \b6_OKctIF[686]  (.D(b4_nUAi[443]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[444]));
    SLE \b6_OKctIF[978]  (.D(b4_nUAi[151]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[152]));
    SLE \b6_OKctIF[1076]  (.D(b4_nUAi[53]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[54]));
    SLE \b6_OKctIF[46]  (.D(b4_nUAi[1083]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1084]));
    SLE \b6_OKctIF[140]  (.D(b4_nUAi[989]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[990]));
    SLE \b6_OKctIF[786]  (.D(b4_nUAi[343]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[344]));
    SLE \b6_OKctIF[487]  (.D(b4_nUAi[642]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[643]));
    SLE \b6_OKctIF[695]  (.D(b4_nUAi[434]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[435]));
    SLE \b6_OKctIF[574]  (.D(b4_nUAi[555]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[556]));
    SLE \b6_OKctIF[967]  (.D(b4_nUAi[162]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[163]));
    SLE \b6_OKctIF[721]  (.D(b4_nUAi[408]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[409]));
    SLE \b6_OKctIF[515]  (.D(b4_nUAi[614]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[615]));
    SLE \b6_OKctIF[864]  (.D(b4_nUAi[265]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[266]));
    SLE \b6_OKctIF[83]  (.D(b4_nUAi[1046]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1047]));
    SLE \b6_OKctIF[385]  (.D(b4_nUAi[744]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[745]));
    SLE \b6_OKctIF[190]  (.D(b4_nUAi[939]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[940]));
    SLE \b6_OKctIF[579]  (.D(b4_nUAi[550]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[551]));
    SLE \b6_OKctIF[82]  (.D(b4_nUAi[1047]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1048]));
    SLE \b6_OKctIF[468]  (.D(b4_nUAi[661]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[662]));
    SLE \b6_OKctIF[224]  (.D(b4_nUAi[905]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[906]));
    SLE \b6_OKctIF[550]  (.D(b4_nUAi[579]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[580]));
    SLE \b6_OKctIF[1119]  (.D(b4_nUAi[10]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[11]));
    SLE \b6_OKctIF[210]  (.D(b4_nUAi[919]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[920]));
    SLE \b6_OKctIF[1018]  (.D(b4_nUAi[111]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[112]));
    SLE \b6_OKctIF[720]  (.D(b4_nUAi[409]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[410]));
    SLE \b6_OKctIF[258]  (.D(b4_nUAi[871]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[872]));
    SLE \b6_OKctIF[916]  (.D(b4_nUAi[213]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[214]));
    SLE \b6_OKctIF[667]  (.D(b4_nUAi[462]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[463]));
    SLE \b6_OKctIF[7]  (.D(b4_nUAi[1122]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1123]));
    SLE \b6_OKctIF[1057]  (.D(b4_nUAi[72]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[73]));
    SLE \b6_OKctIF[540]  (.D(b4_nUAi[589]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[590]));
    SLE \b6_OKctIF[282]  (.D(b4_nUAi[847]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[848]));
    SLE \b6_OKctIF[248]  (.D(b4_nUAi[881]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[882]));
    SLE \b6_OKctIF[922]  (.D(b4_nUAi[207]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[208]));
    SLE \b6_OKctIF[185]  (.D(b4_nUAi[944]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[945]));
    SLE \b6_OKctIF[1085]  (.D(b4_nUAi[44]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[45]));
    SLE \b6_OKctIF[1053]  (.D(b4_nUAi[76]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[77]));
    SLE \b6_OKctIF[586]  (.D(b4_nUAi[543]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[544]));
    SLE \b6_OKctIF[816]  (.D(b4_nUAi[313]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[314]));
    SLE \b6_OKctIF[590]  (.D(b4_nUAi[539]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[540]));
    SLE \b6_OKctIF[373]  (.D(b4_nUAi[756]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[757]));
    SLE \b6_OKctIF[622]  (.D(b4_nUAi[507]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[508]));
    SLE \b6_OKctIF[298]  (.D(b4_nUAi[831]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[832]));
    SLE \b6_OKctIF[531]  (.D(b4_nUAi[598]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[599]));
    SLE \b6_OKctIF[277]  (.D(b4_nUAi[852]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[853]));
    SLE \b6_OKctIF[221]  (.D(b4_nUAi[908]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[909]));
    SLE \b6_OKctIF[624]  (.D(b4_nUAi[505]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[506]));
    SLE \b6_OKctIF[553]  (.D(b4_nUAi[576]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[577]));
    SLE \b6_OKctIF[1091]  (.D(b4_nUAi[38]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[39]));
    SLE \b6_OKctIF[411]  (.D(b4_nUAi[718]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[719]));
    SLE \b6_OKctIF[501]  (.D(b4_nUAi[628]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[629]));
    SLE \b6_OKctIF[129]  (.D(b4_nUAi[1000]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1001]));
    SLE \b6_OKctIF[439]  (.D(b4_nUAi[690]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[691]));
    SLE \b6_OKctIF[452]  (.D(b4_nUAi[677]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[678]));
    SLE \b6_OKctIF[28]  (.D(b4_nUAi[1101]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1102]));
    SLE \b6_OKctIF[650]  (.D(b4_nUAi[479]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[480]));
    SLE \b6_OKctIF[543]  (.D(b4_nUAi[586]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[587]));
    SLE \b6_OKctIF[336]  (.D(b4_nUAi[793]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[794]));
    SLE \b6_OKctIF[6]  (.D(b4_nUAi[1123]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1124]));
    SLE \b6_OKctIF[453]  (.D(b4_nUAi[676]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[677]));
    SLE \b6_OKctIF[768]  (.D(b4_nUAi[361]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[362]));
    SLE \b6_OKctIF[587]  (.D(b4_nUAi[542]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[543]));
    SLE \b6_OKctIF[442]  (.D(b4_nUAi[687]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[688]));
    SLE \b6_OKctIF[184]  (.D(b4_nUAi[945]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[946]));
    SLE \b6_OKctIF[640]  (.D(b4_nUAi[489]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[490]));
    SLE \b6_OKctIF[117]  (.D(b4_nUAi[1012]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1013]));
    SLE \b6_OKctIF[409]  (.D(b4_nUAi[720]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[721]));
    SLE \b6_OKctIF[443]  (.D(b4_nUAi[686]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[687]));
    SLE \b6_OKctIF[593]  (.D(b4_nUAi[536]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[537]));
    SLE \b6_OKctIF[669]  (.D(b4_nUAi[460]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[461]));
    SLE \b6_OKctIF[306]  (.D(b4_nUAi[823]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[824]));
    SLE \b6_OKctIF[259]  (.D(b4_nUAi[870]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[871]));
    SLE \b6_OKctIF[492]  (.D(b4_nUAi[637]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[638]));
    SLE \b6_OKctIF[690]  (.D(b4_nUAi[439]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[440]));
    SLE \b6_OKctIF[493]  (.D(b4_nUAi[636]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[637]));
    SLE \b6_OKctIF[960]  (.D(b4_nUAi[169]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[170]));
    SLE \b6_OKctIF[249]  (.D(b4_nUAi[880]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[881]));
    SLE \b6_OKctIF[1099]  (.D(b4_nUAi[30]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[31]));
    SLE \b6_OKctIF[572]  (.D(b4_nUAi[557]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[558]));
    SLE \b6_OKctIF[934]  (.D(b4_nUAi[195]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[196]));
    SLE \b6_OKctIF[320]  (.D(b4_nUAi[809]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[810]));
    SLE \b6_OKctIF[21]  (.D(b4_nUAi[1108]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1109]));
    SLE \b6_OKctIF[1044]  (.D(b4_nUAi[85]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[86]));
    SLE \b6_OKctIF[1007]  (.D(b4_nUAi[122]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[123]));
    SLE \b6_OKctIF[299]  (.D(b4_nUAi[830]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[831]));
    SLE \b6_OKctIF[861]  (.D(b4_nUAi[268]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[269]));
    SLE \b6_OKctIF[830]  (.D(b4_nUAi[299]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[300]));
    SLE \b6_OKctIF[1003]  (.D(b4_nUAi[126]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[127]));
    SLE \b6_OKctIF[1118]  (.D(b4_nUAi[11]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[12]));
    SLE \b6_OKctIF[1062]  (.D(b4_nUAi[67]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[68]));
    SLE \b6_OKctIF[1050]  (.D(b4_nUAi[79]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[80]));
    SLE \b6_OKctIF[904]  (.D(b4_nUAi[225]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[226]));
    SLE \b6_OKctIF[78]  (.D(b4_nUAi[1051]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1052]));
    SLE \b6_OKctIF[671]  (.D(b4_nUAi[458]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[459]));
    SLE \b6_OKctIF[1066]  (.D(b4_nUAi[63]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[64]));
    SLE \b6_OKctIF[178]  (.D(b4_nUAi[951]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[952]));
    SLE \b6_OKctIF[226]  (.D(b4_nUAi[903]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[904]));
    SLE \b6_OKctIF[800]  (.D(b4_nUAi[329]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[330]));
    SLE \b6_OKctIF[877]  (.D(b4_nUAi[252]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[253]));
    SLE \b6_OKctIF[388]  (.D(b4_nUAi[741]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[742]));
    SLE \b6_OKctIF[152]  (.D(b4_nUAi[977]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[978]));
    SLE \b6_OKctIF[752]  (.D(b4_nUAi[377]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[378]));
    SLE \b6_OKctIF[688]  (.D(b4_nUAi[441]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[442]));
    SLE \b6_OKctIF[424]  (.D(b4_nUAi[705]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[706]));
    SLE \b6_OKctIF[761]  (.D(b4_nUAi[368]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[369]));
    SLE \b6_OKctIF[142]  (.D(b4_nUAi[987]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[988]));
    SLE \b6_OKctIF[476]  (.D(b4_nUAi[653]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[654]));
    SLE \b6_OKctIF[742]  (.D(b4_nUAi[387]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[388]));
    SLE \b6_OKctIF[981]  (.D(b4_nUAi[148]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[149]));
    SLE \b6_OKctIF[3]  (.D(b4_nUAi[1126]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1127]));
    SLE \b6_OKctIF[1015]  (.D(b4_nUAi[114]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[115]));
    SLE \b6_OKctIF[938]  (.D(b4_nUAi[191]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[192]));
    SLE \b6_OKctIF[264]  (.D(b4_nUAi[865]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[866]));
    SLE \b6_OKctIF[192]  (.D(b4_nUAi[937]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[938]));
    SLE \b6_OKctIF[71]  (.D(b4_nUAi[1058]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1059]));
    SLE \b6_OKctIF[792]  (.D(b4_nUAi[337]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[338]));
    SLE \b6_OKctIF[760]  (.D(b4_nUAi[369]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[370]));
    SLE \b6_OKctIF[777]  (.D(b4_nUAi[352]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[353]));
    SLE \b6_OKctIF[121]  (.D(b4_nUAi[1008]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1009]));
    SLE \b6_OKctIF[534]  (.D(b4_nUAi[595]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[596]));
    SLE \b6_OKctIF[683]  (.D(b4_nUAi[446]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[447]));
    SLE \b6_OKctIF[908]  (.D(b4_nUAi[221]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[222]));
    SLE \b6_OKctIF[455]  (.D(b4_nUAi[674]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[675]));
    SLE \b6_OKctIF[962]  (.D(b4_nUAi[167]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[168]));
    SLE \b6_OKctIF[329]  (.D(b4_nUAi[800]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[801]));
    SLE \b6_OKctIF[183]  (.D(b4_nUAi[946]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[947]));
    SLE \b6_OKctIF[852]  (.D(b4_nUAi[277]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[278]));
    SLE \b6_OKctIF[539]  (.D(b4_nUAi[590]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[591]));
    SLE \b6_OKctIF[1107]  (.D(b4_nUAi[22]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[23]));
    SLE \b6_OKctIF[511]  (.D(b4_nUAi[618]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[619]));
    SLE \b6_OKctIF[504]  (.D(b4_nUAi[625]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[626]));
    SLE \b6_OKctIF[445]  (.D(b4_nUAi[684]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[685]));
    SLE \b6_OKctIF[656]  (.D(b4_nUAi[473]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[474]));
    SLE \b6_OKctIF[578]  (.D(b4_nUAi[551]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[552]));
    SLE \b6_OKctIF[8]  (.D(b4_nUAi[1121]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1122]));
    SLE \b6_OKctIF[842]  (.D(b4_nUAi[287]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[288]));
    SLE \b6_OKctIF[662]  (.D(b4_nUAi[467]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[468]));
    SLE \b6_OKctIF[785]  (.D(b4_nUAi[344]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[345]));
    SLE \b6_OKctIF[756]  (.D(b4_nUAi[373]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[374]));
    SLE \b6_OKctIF[457]  (.D(b4_nUAi[672]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[673]));
    SLE \b6_OKctIF[509]  (.D(b4_nUAi[620]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[621]));
    SLE \b6_OKctIF[646]  (.D(b4_nUAi[483]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[484]));
    SLE \b6_OKctIF[495]  (.D(b4_nUAi[634]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[635]));
    SLE \b6_OKctIF[371]  (.D(b4_nUAi[758]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[759]));
    SLE \b6_OKctIF[261]  (.D(b4_nUAi[868]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[869]));
    SLE \b6_OKctIF[664]  (.D(b4_nUAi[465]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[466]));
    SLE \b6_OKctIF[377]  (.D(b4_nUAi[752]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[753]));
    SLE \b6_OKctIF[1000]  (.D(b4_nUAi[129]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[130]));
    SLE \b6_OKctIF[746]  (.D(b4_nUAi[383]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[384]));
    SLE \b6_OKctIF[419]  (.D(b4_nUAi[710]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[711]));
    SLE \b6_OKctIF[892]  (.D(b4_nUAi[237]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[238]));
    SLE \b6_OKctIF[447]  (.D(b4_nUAi[682]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[683]));
    SLE \b6_OKctIF[1129]  (.D(b4_nUAi[0]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1]));
    SLE \b6_OKctIF[1028]  (.D(b4_nUAi[101]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[102]));
    SLE \b6_OKctIF[355]  (.D(b4_nUAi[774]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[775]));
    SLE \b6_OKctIF[316]  (.D(b4_nUAi[813]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[814]));
    SLE \b6_OKctIF[169]  (.D(b4_nUAi[960]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[961]));
    SLE \b6_OKctIF[889]  (.D(b4_nUAi[240]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[241]));
    SLE \b6_OKctIF[1111]  (.D(b4_nUAi[18]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[19]));
    SLE \b6_OKctIF[696]  (.D(b4_nUAi[433]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[434]));
    SLE \b6_OKctIF[26]  (.D(b4_nUAi[1103]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1104]));
    SLE \b6_OKctIF[2]  (.D(b4_nUAi[1127]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1128]));
    SLE \b6_OKctIF[825]  (.D(b4_nUAi[304]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[305]));
    SLE \b6_OKctIF[333]  (.D(b4_nUAi[796]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[797]));
    SLE \b6_OKctIF[989]  (.D(b4_nUAi[140]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[141]));
    SLE \b6_OKctIF[345]  (.D(b4_nUAi[784]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[785]));
    SLE \b6_OKctIF[796]  (.D(b4_nUAi[333]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[334]));
    SLE \b6_OKctIF[497]  (.D(b4_nUAi[632]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[633]));
    SLE \b6_OKctIF[925]  (.D(b4_nUAi[204]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[205]));
    SLE \b6_OKctIF[1041]  (.D(b4_nUAi[88]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[89]));
    SLE \b6_OKctIF[237]  (.D(b4_nUAi[892]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[893]));
    SLE \b6_OKctIF[85]  (.D(b4_nUAi[1044]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1045]));
    SLE \b6_OKctIF[252]  (.D(b4_nUAi[877]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[878]));
    SLE \b6_OKctIF[395]  (.D(b4_nUAi[734]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[735]));
    SLE \b6_OKctIF[303]  (.D(b4_nUAi[826]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[827]));
    SLE \b6_OKctIF[973]  (.D(b4_nUAi[156]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[157]));
    SLE \b6_OKctIF[80]  (.D(b4_nUAi[1049]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1050]));
    SLE \b6_OKctIF[987]  (.D(b4_nUAi[142]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[143]));
    SLE \b6_OKctIF[374]  (.D(b4_nUAi[755]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[756]));
    SLE \b6_OKctIF[155]  (.D(b4_nUAi[974]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[975]));
    SLE \b6_OKctIF[556]  (.D(b4_nUAi[573]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[574]));
    SLE \b6_OKctIF[242]  (.D(b4_nUAi[887]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[888]));
    SLE \b6_OKctIF[884]  (.D(b4_nUAi[245]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[246]));
    SLE \b6_OKctIF[914]  (.D(b4_nUAi[215]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[216]));
    SLE \b6_OKctIF[207]  (.D(b4_nUAi[922]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[923]));
    SLE \b6_OKctIF[145]  (.D(b4_nUAi[984]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[985]));
    SLE \b6_OKctIF[546]  (.D(b4_nUAi[583]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[584]));
    SLE \b6_OKctIF[488]  (.D(b4_nUAi[641]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[642]));
    SLE \b6_OKctIF[360]  (.D(b4_nUAi[769]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[770]));
    SLE \b6_OKctIF[810]  (.D(b4_nUAi[319]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[320]));
    SLE \b6_OKctIF[292]  (.D(b4_nUAi[837]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[838]));
    SLE \b6_OKctIF[687]  (.D(b4_nUAi[442]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[443]));
    SLE \b6_OKctIF[225]  (.D(b4_nUAi[904]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[905]));
    SLE \b6_OKctIF[420]  (.D(b4_nUAi[709]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[710]));
    SLE \b6_OKctIF[195]  (.D(b4_nUAi[934]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[935]));
    SLE \b6_OKctIF[596]  (.D(b4_nUAi[533]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[534]));
    SLE \b6_OKctIF[1049]  (.D(b4_nUAi[80]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[81]));
    SLE \b6_OKctIF[322]  (.D(b4_nUAi[807]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[808]));
    SLE \b6_OKctIF[779]  (.D(b4_nUAi[350]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[351]));
    SLE \b6_OKctIF[76]  (.D(b4_nUAi[1053]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1054]));
    SLE \b6_OKctIF[532]  (.D(b4_nUAi[597]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[598]));
    SLE \b6_OKctIF[266]  (.D(b4_nUAi[863]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[864]));
    SLE \b6_OKctIF[557]  (.D(b4_nUAi[572]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[573]));
    SLE \b6_OKctIF[154]  (.D(b4_nUAi[975]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[976]));
    SLE \b6_OKctIF[464]  (.D(b4_nUAi[665]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[666]));
    SLE \b6_OKctIF[547]  (.D(b4_nUAi[582]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[583]));
    SLE \b6_OKctIF[502]  (.D(b4_nUAi[627]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[628]));
    SLE \b6_OKctIF[144]  (.D(b4_nUAi[985]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[986]));
    SLE \b6_OKctIF[918]  (.D(b4_nUAi[211]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[212]));
    SLE \b6_OKctIF[631]  (.D(b4_nUAi[498]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[499]));
    SLE \b6_OKctIF[138]  (.D(b4_nUAi[991]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[992]));
    SLE \b6_OKctIF[87]  (.D(b4_nUAi[1042]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1043]));
    SLE \b6_OKctIF[873]  (.D(b4_nUAi[256]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[257]));
    SLE \b6_OKctIF[1128]  (.D(b4_nUAi[1]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[2]));
    SLE \b6_OKctIF[597]  (.D(b4_nUAi[532]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[533]));
    SLE \b6_OKctIF[194]  (.D(b4_nUAi[935]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[936]));
    SLE \b6_OKctIF[1104]  (.D(b4_nUAi[25]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[26]));
    SLE \b6_OKctIF[514]  (.D(b4_nUAi[615]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[616]));
    SLE \b6_OKctIF[837]  (.D(b4_nUAi[292]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[293]));
    SLE \b6_OKctIF[1115]  (.D(b4_nUAi[14]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[15]));
    SLE \b6_OKctIF[161]  (.D(b4_nUAi[968]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[969]));
    SLE \b6_OKctIF[788]  (.D(b4_nUAi[341]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[342]));
    SLE \b6_OKctIF[84]  (.D(b4_nUAi[1045]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1046]));
    SLE \b6_OKctIF[1082]  (.D(b4_nUAi[47]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[48]));
    SLE \b6_OKctIF[675]  (.D(b4_nUAi[454]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[455]));
    SLE \b6_OKctIF[601]  (.D(b4_nUAi[528]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[529]));
    SLE \b6_OKctIF[519]  (.D(b4_nUAi[610]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[611]));
    SLE \b6_OKctIF[108]  (.D(b4_nUAi[1021]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1022]));
    SLE \b6_OKctIF[436]  (.D(b4_nUAi[693]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[694]));
    SLE \b6_OKctIF[369]  (.D(b4_nUAi[760]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[761]));
    SLE \b6_OKctIF[807]  (.D(b4_nUAi[322]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[323]));
    SLE \b6_OKctIF[689]  (.D(b4_nUAi[440]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[441]));
    SLE \b6_OKctIF[1086]  (.D(b4_nUAi[43]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[44]));
    SLE \b6_OKctIF[1100]  (.D(b4_nUAi[29]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[30]));
    SLE \b6_OKctIF[170]  (.D(b4_nUAi[959]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[960]));
    SLE \b6_OKctIF[724]  (.D(b4_nUAi[405]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[406]));
    SLE \b6_OKctIF[89]  (.D(b4_nUAi[1040]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1041]));
    SLE \b6_OKctIF[980]  (.D(b4_nUAi[149]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[150]));
    SLE \b6_OKctIF[406]  (.D(b4_nUAi[723]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[724]));
    SLE \b6_OKctIF[358]  (.D(b4_nUAi[771]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[772]));
    SLE \b6_OKctIF[737]  (.D(b4_nUAi[392]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[393]));
    SLE \b6_OKctIF[126]  (.D(b4_nUAi[1003]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1004]));
    SLE \b6_OKctIF[1025]  (.D(b4_nUAi[104]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[105]));
    SLE \b6_OKctIF[658]  (.D(b4_nUAi[471]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[472]));
    SLE \b6_OKctIF[1116]  (.D(b4_nUAi[13]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[14]));
    SLE \b6_OKctIF[348]  (.D(b4_nUAi[781]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[782]));
    SLE \b6_OKctIF[648]  (.D(b4_nUAi[481]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[482]));
    SLE \b6_OKctIF[881]  (.D(b4_nUAi[248]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[249]));
    SLE \b6_OKctIF[313]  (.D(b4_nUAi[816]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[817]));
    SLE \b6_OKctIF[951]  (.D(b4_nUAi[178]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[179]));
    SLE \b6_OKctIF[63]  (.D(b4_nUAi[1066]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1067]));
    SLE \b6_OKctIF[1037]  (.D(b4_nUAi[92]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[93]));
    SLE \b6_OKctIF[707]  (.D(b4_nUAi[422]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[423]));
    SLE \b6_OKctIF[723]  (.D(b4_nUAi[406]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[407]));
    SLE \b6_OKctIF[865]  (.D(b4_nUAi[264]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[265]));
    SLE \b6_OKctIF[538]  (.D(b4_nUAi[591]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[592]));
    SLE \b6_OKctIF[62]  (.D(b4_nUAi[1067]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1068]));
    SLE \b6_OKctIF[398]  (.D(b4_nUAi[731]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[732]));
    SLE \b6_OKctIF[1033]  (.D(b4_nUAi[96]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[97]));
    SLE \b6_OKctIF[941]  (.D(b4_nUAi[188]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[189]));
    SLE \b6_OKctIF[570]  (.D(b4_nUAi[559]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[560]));
    SLE \b6_OKctIF[965]  (.D(b4_nUAi[164]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[165]));
    SLE \b6_OKctIF[828]  (.D(b4_nUAi[301]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[302]));
    SLE \b6_OKctIF[217]  (.D(b4_nUAi[912]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[913]));
    SLE \b6_OKctIF[1]  (.D(b4_nUAi[1128]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1129]));
    SLE \b6_OKctIF[698]  (.D(b4_nUAi[431]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[432]));
    SLE \b6_OKctIF[223]  (.D(b4_nUAi[906]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[907]));
    SLE \b6_OKctIF[278]  (.D(b4_nUAi[851]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[852]));
    SLE \b6_OKctIF[331]  (.D(b4_nUAi[798]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[799]));
    SLE \b6_OKctIF[653]  (.D(b4_nUAi[476]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[477]));
    SLE \b6_OKctIF[337]  (.D(b4_nUAi[792]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[793]));
    SLE \b6_OKctIF[1098]  (.D(b4_nUAi[31]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[32]));
    SLE \b6_OKctIF[508]  (.D(b4_nUAi[621]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[622]));
    SLE \b6_OKctIF[991]  (.D(b4_nUAi[138]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[139]));
    SLE \b6_OKctIF[781]  (.D(b4_nUAi[348]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[349]));
    SLE \b6_OKctIF[153]  (.D(b4_nUAi[976]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[977]));
    SLE \b6_OKctIF[643]  (.D(b4_nUAi[486]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[487]));
    SLE \b6_OKctIF[1077]  (.D(b4_nUAi[52]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[53]));
    SLE \b6_OKctIF[525]  (.D(b4_nUAi[604]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[605]));
    SLE \b6_OKctIF[301]  (.D(b4_nUAi[828]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[829]));
    SLE \b6_OKctIF[307]  (.D(b4_nUAi[822]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[823]));
    SLE \b6_OKctIF[143]  (.D(b4_nUAi[986]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[987]));
    SLE \b6_OKctIF[755]  (.D(b4_nUAi[374]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[375]));
    SLE \b6_OKctIF[1073]  (.D(b4_nUAi[56]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[57]));
    SLE \b6_OKctIF[1121]  (.D(b4_nUAi[8]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[9]));
    SLE \b6_OKctIF[284]  (.D(b4_nUAi[845]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[846]));
    SLE \b6_OKctIF[693]  (.D(b4_nUAi[436]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[437]));
    SLE \b6_OKctIF[1054]  (.D(b4_nUAi[75]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[76]));
    SLE \b6_OKctIF[780]  (.D(b4_nUAi[349]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[350]));
    SLE \b6_OKctIF[745]  (.D(b4_nUAi[384]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[385]));
    SLE \b6_OKctIF[265]  (.D(b4_nUAi[864]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[865]));
    SLE \b6_OKctIF[460]  (.D(b4_nUAi[669]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[670]));
    SLE \b6_OKctIF[933]  (.D(b4_nUAi[196]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[197]));
    SLE \b6_OKctIF[573]  (.D(b4_nUAi[556]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[557]));
    SLE \b6_OKctIF[193]  (.D(b4_nUAi[936]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[937]));
    SLE \b6_OKctIF[13]  (.D(b4_nUAi[1116]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1117]));
    SLE \b6_OKctIF[362]  (.D(b4_nUAi[767]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[768]));
    SLE \b6_OKctIF[334]  (.D(b4_nUAi[795]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[796]));
    SLE \b6_OKctIF[220]  (.D(b4_nUAi[909]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[910]));
    SLE \b6_OKctIF[512]  (.D(b4_nUAi[617]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[618]));
    SLE \b6_OKctIF[926]  (.D(b4_nUAi[203]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[204]));
    SLE \b6_OKctIF[859]  (.D(b4_nUAi[270]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[271]));
    SLE \b6_OKctIF[472]  (.D(b4_nUAi[657]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[658]));
    SLE \b6_OKctIF[982]  (.D(b4_nUAi[147]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[148]));
    SLE \b6_OKctIF[12]  (.D(b4_nUAi[1117]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1118]));
    SLE \b6_OKctIF[670]  (.D(b4_nUAi[459]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[460]));
    SLE \b6_OKctIF[795]  (.D(b4_nUAi[334]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[335]));
    SLE \b6_OKctIF[959]  (.D(b4_nUAi[170]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[171]));
    SLE \b6_OKctIF[473]  (.D(b4_nUAi[656]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[657]));
    SLE \b6_OKctIF[903]  (.D(b4_nUAi[226]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[227]));
    SLE \b6_OKctIF[849]  (.D(b4_nUAi[280]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[281]));
    SLE \b6_OKctIF[304]  (.D(b4_nUAi[825]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[826]));
    SLE \b6_OKctIF[682]  (.D(b4_nUAi[447]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[448]));
    SLE \b6_OKctIF[949]  (.D(b4_nUAi[180]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[181]));
    SLE \b6_OKctIF[826]  (.D(b4_nUAi[303]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[304]));
    SLE \b6_OKctIF[279]  (.D(b4_nUAi[850]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[851]));
    SLE \b6_OKctIF[899]  (.D(b4_nUAi[230]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[231]));
    SLE \b6_OKctIF[1012]  (.D(b4_nUAi[117]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[118]));
    SLE \b6_OKctIF[957]  (.D(b4_nUAi[172]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[173]));
    SLE \b6_OKctIF[611]  (.D(b4_nUAi[518]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[519]));
    SLE \b6_OKctIF[281]  (.D(b4_nUAi[848]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[849]));
    SLE \b6_OKctIF[93]  (.D(b4_nUAi[1036]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1037]));
    SLE \b6_OKctIF[118]  (.D(b4_nUAi[1011]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1012]));
    SLE \b6_OKctIF[739]  (.D(b4_nUAi[390]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[391]));
    SLE \b6_OKctIF[684]  (.D(b4_nUAi[445]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[446]));
    SLE \b6_OKctIF[999]  (.D(b4_nUAi[130]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[131]));
    SLE \b6_OKctIF[854]  (.D(b4_nUAi[275]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[276]));
    SLE \b6_OKctIF[817]  (.D(b4_nUAi[312]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[313]));
    SLE \b6_OKctIF[1016]  (.D(b4_nUAi[113]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[114]));
    SLE \b6_OKctIF[92]  (.D(b4_nUAi[1037]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1038]));
    SLE \b6_OKctIF[189]  (.D(b4_nUAi[940]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[941]));
    SLE \b6_OKctIF[947]  (.D(b4_nUAi[182]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[183]));
    SLE \b6_OKctIF[1030]  (.D(b4_nUAi[99]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[100]));
    SLE \b6_OKctIF[421]  (.D(b4_nUAi[708]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[709]));
    SLE \b6_OKctIF[458]  (.D(b4_nUAi[671]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[672]));
    SLE \b6_OKctIF[844]  (.D(b4_nUAi[285]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[286]));
    SLE \b6_OKctIF[709]  (.D(b4_nUAi[420]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[421]));
    SLE \b6_OKctIF[1103]  (.D(b4_nUAi[26]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[27]));
    SLE \b6_OKctIF[416]  (.D(b4_nUAi[713]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[714]));
    SLE \b6_OKctIF[997]  (.D(b4_nUAi[132]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[133]));
    SLE \b6_OKctIF[448]  (.D(b4_nUAi[681]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[682]));
    SLE \b6_OKctIF[657]  (.D(b4_nUAi[472]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[473]));
    SLE \b6_OKctIF[127]  (.D(b4_nUAi[1002]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1003]));
    SLE \b6_OKctIF[894]  (.D(b4_nUAi[235]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[236]));
    SLE \b6_OKctIF[764]  (.D(b4_nUAi[365]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[366]));
    SLE \b6_OKctIF[647]  (.D(b4_nUAi[482]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[483]));
    SLE \b6_OKctIF[833]  (.D(b4_nUAi[296]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[297]));
    SLE \b6_OKctIF[717]  (.D(b4_nUAi[412]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[413]));
    SLE \b6_OKctIF[498]  (.D(b4_nUAi[631]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[632]));
    SLE \b6_OKctIF[1070]  (.D(b4_nUAi[59]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[60]));
    SLE \b6_OKctIF[172]  (.D(b4_nUAi[957]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[958]));
    SLE \b6_OKctIF[166]  (.D(b4_nUAi[963]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[964]));
    SLE \b6_OKctIF[1004]  (.D(b4_nUAi[125]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[126]));
    SLE \b6_OKctIF[772]  (.D(b4_nUAi[357]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[358]));
    SLE \b6_OKctIF[697]  (.D(b4_nUAi[432]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[433]));
    SLE \b6_OKctIF[380]  (.D(b4_nUAi[749]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[750]));
    SLE \b6_OKctIF[635]  (.D(b4_nUAi[494]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[495]));
    SLE \b6_OKctIF[803]  (.D(b4_nUAi[326]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[327]));
    SLE \b6_OKctIF[1102]  (.D(b4_nUAi[27]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[28]));
    SLE \b6_OKctIF[1125]  (.D(b4_nUAi[4]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[5]));
    SLE \b6_OKctIF[518]  (.D(b4_nUAi[611]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[612]));
    SLE \b6_OKctIF[130]  (.D(b4_nUAi[999]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1000]));
    SLE \b6_OKctIF[763]  (.D(b4_nUAi[366]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[367]));
    SLE \b6_OKctIF[605]  (.D(b4_nUAi[524]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[525]));
    SLE \b6_OKctIF[868]  (.D(b4_nUAi[261]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[262]));
    SLE \b6_OKctIF[311]  (.D(b4_nUAi[818]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[819]));
    SLE \b6_OKctIF[263]  (.D(b4_nUAi[866]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[867]));
    SLE \b6_OKctIF[1095]  (.D(b4_nUAi[34]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[35]));
    SLE \b6_OKctIF[317]  (.D(b4_nUAi[812]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[813]));
    SLE \b6_OKctIF[286]  (.D(b4_nUAi[843]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[844]));
    SLE \b6_OKctIF[100]  (.D(b4_nUAi[1029]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1030]));
    SLE \b6_OKctIF[758]  (.D(b4_nUAi[371]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[372]));
    SLE \b6_OKctIF[1051]  (.D(b4_nUAi[78]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[79]));
    SLE \b6_OKctIF[484]  (.D(b4_nUAi[645]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[646]));
    SLE \b6_OKctIF[475]  (.D(b4_nUAi[654]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[655]));
    SLE \b6_OKctIF[33]  (.D(b4_nUAi[1096]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1097]));
    SLE \b6_OKctIF[1067]  (.D(b4_nUAi[62]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[63]));
    SLE \b6_OKctIF[872]  (.D(b4_nUAi[257]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[258]));
    SLE \b6_OKctIF[748]  (.D(b4_nUAi[381]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[382]));
    SLE \b6_OKctIF[659]  (.D(b4_nUAi[470]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[471]));
    SLE \b6_OKctIF[32]  (.D(b4_nUAi[1097]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1098]));
    SLE \b6_OKctIF[565]  (.D(b4_nUAi[564]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[565]));
    SLE \b6_OKctIF[1126]  (.D(b4_nUAi[3]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[4]));
    SLE \b6_OKctIF[1063]  (.D(b4_nUAi[66]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[67]));
    SLE \b6_OKctIF[676]  (.D(b4_nUAi[453]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[454]));
    SLE \b6_OKctIF[649]  (.D(b4_nUAi[480]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[481]));
    SLE \b6_OKctIF[530]  (.D(b4_nUAi[599]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[600]));
    SLE \b6_OKctIF[950]  (.D(b4_nUAi[179]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[180]));
    SLE \b6_OKctIF[776]  (.D(b4_nUAi[353]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[354]));
    SLE \b6_OKctIF[1048]  (.D(b4_nUAi[81]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[82]));
    SLE \b6_OKctIF[798]  (.D(b4_nUAi[331]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[332]));
    SLE \b6_OKctIF[477]  (.D(b4_nUAi[652]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[653]));
    SLE \b6_OKctIF[238]  (.D(b4_nUAi[891]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[892]));
    SLE \b6_OKctIF[913]  (.D(b4_nUAi[216]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[217]));
    SLE \b6_OKctIF[314]  (.D(b4_nUAi[815]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[816]));
    SLE \b6_OKctIF[940]  (.D(b4_nUAi[189]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[190]));
    SLE \b6_OKctIF[181]  (.D(b4_nUAi[948]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[949]));
    SLE \b6_OKctIF[699]  (.D(b4_nUAi[430]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[431]));
    SLE \b6_OKctIF[500]  (.D(b4_nUAi[629]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[630]));
    SLE \b6_OKctIF[260]  (.D(b4_nUAi[869]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[870]));
    SLE \b6_OKctIF[375]  (.D(b4_nUAi[754]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[755]));
    SLE \b6_OKctIF[966]  (.D(b4_nUAi[163]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[164]));
    SLE \b6_OKctIF[851]  (.D(b4_nUAi[278]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[279]));
    SLE \b6_OKctIF[208]  (.D(b4_nUAi[921]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[922]));
    SLE \b6_OKctIF[1059]  (.D(b4_nUAi[70]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[71]));
    SLE \b6_OKctIF[389]  (.D(b4_nUAi[740]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[741]));
    SLE \b6_OKctIF[990]  (.D(b4_nUAi[139]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[140]));
    SLE \b6_OKctIF[841]  (.D(b4_nUAi[288]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[289]));
    SLE \b6_OKctIF[1130]  (.D(b4_PLyF), .CLK(IICE_comm2iice[11]), .EN(
        b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[0]));
    SLE \b6_OKctIF[866]  (.D(b4_nUAi[263]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[264]));
    SLE \b6_OKctIF[521]  (.D(b4_nUAi[608]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[609]));
    SLE \b6_OKctIF[719]  (.D(b4_nUAi[410]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[411]));
    SLE \b6_OKctIF[272]  (.D(b4_nUAi[857]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[858]));
    SLE \b6_OKctIF[533]  (.D(b4_nUAi[596]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[597]));
    SLE \b6_OKctIF[891]  (.D(b4_nUAi[238]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[239]));
    SLE \b6_OKctIF[65]  (.D(b4_nUAi[1064]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1065]));
    SLE \b6_OKctIF[751]  (.D(b4_nUAi[378]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[379]));
    SLE \b6_OKctIF[60]  (.D(b4_nUAi[1069]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1070]));
    SLE \b6_OKctIF[175]  (.D(b4_nUAi[954]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[955]));
    SLE \b6_OKctIF[576]  (.D(b4_nUAi[553]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[554]));
    SLE \b6_OKctIF[432]  (.D(b4_nUAi[697]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[698]));
    SLE \b6_OKctIF[630]  (.D(b4_nUAi[499]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[500]));
    SLE \b6_OKctIF[741]  (.D(b4_nUAi[388]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[389]));
    SLE \b6_OKctIF[429]  (.D(b4_nUAi[700]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[701]));
    SLE \b6_OKctIF[433]  (.D(b4_nUAi[696]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[697]));
    SLE \b6_OKctIF[461]  (.D(b4_nUAi[668]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[669]));
    SLE \b6_OKctIF[503]  (.D(b4_nUAi[626]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[627]));
    SLE \b6_OKctIF[326]  (.D(b4_nUAi[803]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[804]));
    SLE \b6_OKctIF[885]  (.D(b4_nUAi[244]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[245]));
    SLE \b6_OKctIF[254]  (.D(b4_nUAi[875]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[876]));
    SLE \b6_OKctIF[1001]  (.D(b4_nUAi[128]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[129]));
    SLE \b6_OKctIF[985]  (.D(b4_nUAi[144]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[145]));
    SLE \b6_OKctIF[402]  (.D(b4_nUAi[727]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[728]));
    SLE \b6_OKctIF[600]  (.D(b4_nUAi[529]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[530]));
    SLE \b6_OKctIF[750]  (.D(b4_nUAi[379]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[380]));
    SLE \b6_OKctIF[791]  (.D(b4_nUAi[338]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[339]));
    SLE \b6_OKctIF[403]  (.D(b4_nUAi[726]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[727]));
    SLE \b6_OKctIF[239]  (.D(b4_nUAi[890]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[891]));
    SLE \b6_OKctIF[244]  (.D(b4_nUAi[885]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[886]));
    SLE \b6_OKctIF[167]  (.D(b4_nUAi[962]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[963]));
    SLE \b6_OKctIF[88]  (.D(b4_nUAi[1041]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1042]));
    SLE \b6_OKctIF[813]  (.D(b4_nUAi[316]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[317]));
    SLE \b6_OKctIF[740]  (.D(b4_nUAi[389]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[390]));
    SLE \b6_OKctIF[952]  (.D(b4_nUAi[177]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[178]));
    SLE \b6_OKctIF[1060]  (.D(b4_nUAi[69]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[70]));
    SLE \b6_OKctIF[1022]  (.D(b4_nUAi[107]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[108]));
    SLE \b6_OKctIF[294]  (.D(b4_nUAi[835]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[836]));
    SLE \b6_OKctIF[209]  (.D(b4_nUAi[920]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[921]));
    SLE \b6_OKctIF[577]  (.D(b4_nUAi[552]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[553]));
    SLE \b6_OKctIF[942]  (.D(b4_nUAi[187]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[188]));
    SLE \b6_OKctIF[615]  (.D(b4_nUAi[514]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[515]));
    SLE \b6_OKctIF[174]  (.D(b4_nUAi[955]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[956]));
    SLE \b6_OKctIF[790]  (.D(b4_nUAi[339]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[340]));
    SLE \b6_OKctIF[652]  (.D(b4_nUAi[477]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[478]));
    SLE \b6_OKctIF[1026]  (.D(b4_nUAi[103]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[104]));
    SLE \b6_OKctIF[924]  (.D(b4_nUAi[205]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[206]));
    SLE \b6_OKctIF[15]  (.D(b4_nUAi[1114]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1115]));
    SLE \b6_OKctIF[4]  (.D(b4_nUAi[1125]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1126]));
    SLE \b6_OKctIF[10]  (.D(b4_nUAi[1119]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1120]));
    SLE \b6_OKctIF[110]  (.D(b4_nUAi[1019]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1020]));
    SLE \b6_OKctIF[642]  (.D(b4_nUAi[487]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[488]));
    SLE \b6_OKctIF[1009]  (.D(b4_nUAi[120]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[121]));
    SLE \b6_OKctIF[251]  (.D(b4_nUAi[878]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[879]));
    SLE \b6_OKctIF[992]  (.D(b4_nUAi[137]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[138]));
    SLE \b6_OKctIF[285]  (.D(b4_nUAi[844]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[845]));
    SLE \b6_OKctIF[820]  (.D(b4_nUAi[309]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[310]));
    SLE \b6_OKctIF[654]  (.D(b4_nUAi[475]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[476]));
    SLE \b6_OKctIF[480]  (.D(b4_nUAi[649]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[650]));
    SLE \b6_OKctIF[382]  (.D(b4_nUAi[747]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[748]));
    SLE \b6_OKctIF[159]  (.D(b4_nUAi[970]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[971]));
    SLE \b6_OKctIF[241]  (.D(b4_nUAi[888]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[889]));
    SLE \b6_OKctIF[81]  (.D(b4_nUAi[1048]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1049]));
    SLE \b6_OKctIF[67]  (.D(b4_nUAi[1062]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1063]));
    SLE \b6_OKctIF[644]  (.D(b4_nUAi[485]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[486]));
    SLE \b6_OKctIF[692]  (.D(b4_nUAi[437]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[438]));
    SLE \b6_OKctIF[132]  (.D(b4_nUAi[997]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[998]));
    SLE \b6_OKctIF[149]  (.D(b4_nUAi[980]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[981]));
    SLE \b6_OKctIF[732]  (.D(b4_nUAi[397]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[398]));
    SLE \b6_OKctIF[95]  (.D(b4_nUAi[1034]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1035]));
    SLE \b6_OKctIF[64]  (.D(b4_nUAi[1065]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1066]));
    SLE \b6_OKctIF[291]  (.D(b4_nUAi[838]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[839]));
    SLE \b6_OKctIF[694]  (.D(b4_nUAi[435]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[436]));
    SLE \b6_OKctIF[90]  (.D(b4_nUAi[1039]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1040]));
    SLE \b6_OKctIF[102]  (.D(b4_nUAi[1027]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1028]));
    SLE \b6_OKctIF[199]  (.D(b4_nUAi[930]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[931]));
    SLE \b6_OKctIF[510]  (.D(b4_nUAi[619]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[620]));
    SLE \b6_OKctIF[702]  (.D(b4_nUAi[427]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[428]));
    SLE \b6_OKctIF[1045]  (.D(b4_nUAi[84]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[85]));
    SLE \b6_OKctIF[218]  (.D(b4_nUAi[911]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[912]));
    SLE \b6_OKctIF[69]  (.D(b4_nUAi[1060]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1061]));
    SLE \b6_OKctIF[928]  (.D(b4_nUAi[201]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[202]));
    SLE \b6_OKctIF[378]  (.D(b4_nUAi[751]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[752]));
    SLE \b6_OKctIF[678]  (.D(b4_nUAi[451]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[452]));
    SLE \b6_OKctIF[350]  (.D(b4_nUAi[779]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[780]));
    SLE \b6_OKctIF[524]  (.D(b4_nUAi[605]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[606]));
    SLE \b6_OKctIF[435]  (.D(b4_nUAi[694]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[695]));
    SLE \b6_OKctIF[832]  (.D(b4_nUAi[297]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[298]));
    SLE \b6_OKctIF[971]  (.D(b4_nUAi[158]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[159]));
    SLE \b6_OKctIF[340]  (.D(b4_nUAi[789]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[790]));
    SLE \b6_OKctIF[17]  (.D(b4_nUAi[1112]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1113]));
    SLE \b6_OKctIF[529]  (.D(b4_nUAi[600]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[601]));
    SLE \b6_OKctIF[636]  (.D(b4_nUAi[493]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[494]));
    SLE \b6_OKctIF[784]  (.D(b4_nUAi[345]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[346]));
    SLE \b6_OKctIF[405]  (.D(b4_nUAi[724]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[725]));
    SLE \b6_OKctIF[736]  (.D(b4_nUAi[393]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[394]));
    SLE \b6_OKctIF[437]  (.D(b4_nUAi[692]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[693]));
    SLE \b6_OKctIF[802]  (.D(b4_nUAi[327]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[328]));
    SLE \b6_OKctIF[390]  (.D(b4_nUAi[739]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[740]));
    SLE \b6_OKctIF[256]  (.D(b4_nUAi[873]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[874]));
    SLE \b6_OKctIF[561]  (.D(b4_nUAi[568]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[569]));
    SLE \b6_OKctIF[513]  (.D(b4_nUAi[616]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[617]));
    SLE \b6_OKctIF[14]  (.D(b4_nUAi[1115]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1116]));
    SLE \b6_OKctIF[673]  (.D(b4_nUAi[456]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[457]));
    SLE \b6_OKctIF[186]  (.D(b4_nUAi[943]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[944]));
    SLE \b6_OKctIF[1087]  (.D(b4_nUAi[42]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[43]));
    SLE \b6_OKctIF[606]  (.D(b4_nUAi[523]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[524]));
    SLE \b6_OKctIF[412]  (.D(b4_nUAi[717]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[718]));
    SLE \b6_OKctIF[454]  (.D(b4_nUAi[675]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[676]));
    SLE \b6_OKctIF[246]  (.D(b4_nUAi[883]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[884]));
    SLE \b6_OKctIF[610]  (.D(b4_nUAi[519]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[520]));
    SLE \b6_OKctIF[335]  (.D(b4_nUAi[794]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[795]));
    SLE \b6_OKctIF[173]  (.D(b4_nUAi[956]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[957]));
    SLE \b6_OKctIF[706]  (.D(b4_nUAi[423]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[424]));
    SLE \b6_OKctIF[1083]  (.D(b4_nUAi[46]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[47]));
    SLE \b6_OKctIF[1034]  (.D(b4_nUAi[95]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[96]));
    SLE \b6_OKctIF[413]  (.D(b4_nUAi[716]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[717]));
    SLE \b6_OKctIF[407]  (.D(b4_nUAi[722]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[723]));
    SLE \b6_OKctIF[19]  (.D(b4_nUAi[1110]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1111]));
    SLE \b6_OKctIF[444]  (.D(b4_nUAi[685]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[686]));
    SLE \b6_OKctIF[469]  (.D(b4_nUAi[660]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[661]));
    SLE \b6_OKctIF[97]  (.D(b4_nUAi[1032]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1033]));
    SLE \b6_OKctIF[783]  (.D(b4_nUAi[346]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[347]));
    SLE \b6_OKctIF[775]  (.D(b4_nUAi[354]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[355]));
    SLE \b6_OKctIF[366]  (.D(b4_nUAi[763]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[764]));
    SLE \b6_OKctIF[296]  (.D(b4_nUAi[833]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[834]));
    SLE \b6_OKctIF[323]  (.D(b4_nUAi[806]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[807]));
    SLE \b6_OKctIF[305]  (.D(b4_nUAi[824]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[825]));
    SLE \b6_OKctIF[219]  (.D(b4_nUAi[910]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[911]));
    SLE \b6_OKctIF[888]  (.D(b4_nUAi[241]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[242]));
    SLE \b6_OKctIF[35]  (.D(b4_nUAi[1094]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1095]));
    SLE \b6_OKctIF[283]  (.D(b4_nUAi[846]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[847]));
    SLE \b6_OKctIF[94]  (.D(b4_nUAi[1035]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1036]));
    SLE \b6_OKctIF[494]  (.D(b4_nUAi[635]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[636]));
    SLE \b6_OKctIF[232]  (.D(b4_nUAi[897]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[898]));
    SLE \b6_OKctIF[30]  (.D(b4_nUAi[1099]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1100]));
    SLE \b6_OKctIF[151]  (.D(b4_nUAi[978]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[979]));
    SLE \b6_OKctIF[227]  (.D(b4_nUAi[902]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[903]));
    SLE \b6_OKctIF[135]  (.D(b4_nUAi[994]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[995]));
    SLE \b6_OKctIF[879]  (.D(b4_nUAi[250]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[251]));
    SLE \b6_OKctIF[86]  (.D(b4_nUAi[1043]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1044]));
    SLE \b6_OKctIF[536]  (.D(b4_nUAi[593]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[594]));
    SLE \b6_OKctIF[1074]  (.D(b4_nUAi[55]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[56]));
    SLE \b6_OKctIF[141]  (.D(b4_nUAi[988]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[989]));
    SLE \b6_OKctIF[359]  (.D(b4_nUAi[770]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[771]));
    SLE \b6_OKctIF[99]  (.D(b4_nUAi[1030]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1031]));
    SLE \b6_OKctIF[979]  (.D(b4_nUAi[150]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[151]));
    SLE \b6_OKctIF[202]  (.D(b4_nUAi[927]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[928]));
    SLE \b6_OKctIF[585]  (.D(b4_nUAi[544]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[545]));
    SLE \b6_OKctIF[349]  (.D(b4_nUAi[780]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[781]));
    SLE \b6_OKctIF[105]  (.D(b4_nUAi[1024]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1025]));
    SLE \b6_OKctIF[506]  (.D(b4_nUAi[623]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[624]));
    SLE \b6_OKctIF[964]  (.D(b4_nUAi[165]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[166]));
    SLE \b6_OKctIF[191]  (.D(b4_nUAi[938]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[939]));
    SLE \b6_OKctIF[977]  (.D(b4_nUAi[152]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[153]));
    SLE \b6_OKctIF[860]  (.D(b4_nUAi[269]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[270]));
    SLE \b6_OKctIF[399]  (.D(b4_nUAi[730]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[731]));
    SLE \b6_OKctIF[874]  (.D(b4_nUAi[255]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[256]));
    SLE \b6_OKctIF[280]  (.D(b4_nUAi[849]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[850]));
    SLE \b6_OKctIF[53]  (.D(b4_nUAi[1076]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1077]));
    SLE \b6_OKctIF[1092]  (.D(b4_nUAi[37]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[38]));
    SLE \b6_OKctIF[986]  (.D(b4_nUAi[143]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[144]));
    SLE \b6_OKctIF[112]  (.D(b4_nUAi[1017]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1018]));
    SLE \b6_OKctIF[712]  (.D(b4_nUAi[417]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[418]));
    SLE \b6_OKctIF[537]  (.D(b4_nUAi[592]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[593]));
    SLE \b6_OKctIF[52]  (.D(b4_nUAi[1077]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1078]));
    SLE \b6_OKctIF[522]  (.D(b4_nUAi[607]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[608]));
    SLE \b6_OKctIF[478]  (.D(b4_nUAi[651]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[652]));
    SLE \b6_OKctIF[855]  (.D(b4_nUAi[274]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[275]));
    SLE \b6_OKctIF[134]  (.D(b4_nUAi[995]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[996]));
    SLE \b6_OKctIF[1096]  (.D(b4_nUAi[33]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[34]));
    SLE \b6_OKctIF[955]  (.D(b4_nUAi[174]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[175]));
    SLE \b6_OKctIF[845]  (.D(b4_nUAi[284]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[285]));
    SLE \b6_OKctIF[677]  (.D(b4_nUAi[452]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[453]));
    SLE \b6_OKctIF[886]  (.D(b4_nUAi[243]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[244]));
    SLE \b6_OKctIF[945]  (.D(b4_nUAi[184]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[185]));
    SLE \b6_OKctIF[507]  (.D(b4_nUAi[622]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[623]));
    SLE \b6_OKctIF[1080]  (.D(b4_nUAi[49]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[50]));
    SLE \b6_OKctIF[104]  (.D(b4_nUAi[1025]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1026]));
    SLE \b6_OKctIF[37]  (.D(b4_nUAi[1092]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1093]));
    SLE \b6_OKctIF[895]  (.D(b4_nUAi[234]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[235]));
    SLE \b6_OKctIF[621]  (.D(b4_nUAi[508]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[509]));
    SLE \b6_OKctIF[128]  (.D(b4_nUAi[1001]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1002]));
    SLE \b6_OKctIF[968]  (.D(b4_nUAi[161]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[162]));
    SLE \b6_OKctIF[995]  (.D(b4_nUAi[134]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[135]));
    SLE \b6_OKctIF[481]  (.D(b4_nUAi[648]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[649]));
    SLE \b6_OKctIF[415]  (.D(b4_nUAi[714]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[715]));
    SLE \b6_OKctIF[34]  (.D(b4_nUAi[1095]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1096]));
    SLE \b6_OKctIF[827]  (.D(b4_nUAi[302]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[303]));
    SLE \b6_OKctIF[1058]  (.D(b4_nUAi[71]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[72]));
    SLE \b6_OKctIF[812]  (.D(b4_nUAi[317]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[318]));
    SLE \b6_OKctIF[564]  (.D(b4_nUAi[565]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[566]));
    SLE \b6_OKctIF[1017]  (.D(b4_nUAi[112]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[113]));
    SLE \b6_OKctIF[616]  (.D(b4_nUAi[513]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[514]));
    SLE \b6_OKctIF[255]  (.D(b4_nUAi[874]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[875]));
    SLE \b6_OKctIF[450]  (.D(b4_nUAi[679]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[680]));
    SLE \b6_OKctIF[426]  (.D(b4_nUAi[703]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[704]));
    SLE \b6_OKctIF[39]  (.D(b4_nUAi[1090]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1091]));
    SLE \b6_OKctIF[1031]  (.D(b4_nUAi[98]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[99]));
    SLE \b6_OKctIF[352]  (.D(b4_nUAi[777]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[778]));
    SLE \b6_OKctIF[187]  (.D(b4_nUAi[942]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[943]));
    SLE \b6_OKctIF[569]  (.D(b4_nUAi[560]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[561]));
    SLE \b6_OKctIF[716]  (.D(b4_nUAi[413]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[414]));
    SLE \b6_OKctIF[1013]  (.D(b4_nUAi[116]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[117]));
    SLE \b6_OKctIF[417]  (.D(b4_nUAi[712]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[713]));
    SLE \b6_OKctIF[245]  (.D(b4_nUAi[884]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[885]));
    SLE \b6_OKctIF[440]  (.D(b4_nUAi[689]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[690]));
    SLE \b6_OKctIF[342]  (.D(b4_nUAi[787]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[788]));
    SLE \b6_OKctIF[338]  (.D(b4_nUAi[791]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[792]));
    SLE \b6_OKctIF[638]  (.D(b4_nUAi[491]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[492]));
    SLE \b6_OKctIF[778]  (.D(b4_nUAi[351]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[352]));
    SLE \b6_OKctIF[43]  (.D(b4_nUAi[1086]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1087]));
    SLE \b6_OKctIF[315]  (.D(b4_nUAi[814]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[815]));
    SLE \b6_OKctIF[727]  (.D(b4_nUAi[402]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[403]));
    SLE \b6_OKctIF[295]  (.D(b4_nUAi[834]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[835]));
    SLE \b6_OKctIF[490]  (.D(b4_nUAi[639]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[640]));
    SLE \b6_OKctIF[42]  (.D(b4_nUAi[1087]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1088]));
    SLE \b6_OKctIF[679]  (.D(b4_nUAi[450]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[451]));
    SLE \b6_OKctIF[392]  (.D(b4_nUAi[737]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[738]));
    SLE \b6_OKctIF[931]  (.D(b4_nUAi[198]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[199]));
    SLE \b6_OKctIF[308]  (.D(b4_nUAi[821]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[822]));
    SLE \b6_OKctIF[608]  (.D(b4_nUAi[521]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[522]));
    SLE \b6_OKctIF[1071]  (.D(b4_nUAi[58]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[59]));
    CFG2 #( .INIT(4'h8) )  b6_OKctIF4 (.A(b8_PSyiBgYG), .B(
        IICE_comm2iice[10]), .Y(b6_OKctIF4_net_1));
    SLE \b6_OKctIF[970]  (.D(b4_nUAi[159]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[160]));
    SLE \b6_OKctIF[363]  (.D(b4_nUAi[766]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[767]));
    SLE \b6_OKctIF[1039]  (.D(b4_nUAi[90]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[91]));
    SLE \b6_OKctIF[528]  (.D(b4_nUAi[601]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[602]));
    SLE \b6_OKctIF[212]  (.D(b4_nUAi[917]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[918]));
    SLE \b6_OKctIF[901]  (.D(b4_nUAi[228]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[229]));
    SLE \b6_OKctIF[633]  (.D(b4_nUAi[496]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[497]));
    SLE \b6_OKctIF[115]  (.D(b4_nUAi[1014]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1015]));
    SLE \b6_OKctIF[516]  (.D(b4_nUAi[613]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[614]));
    SLE \b6_OKctIF[267]  (.D(b4_nUAi[862]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[863]));
    SLE \b6_OKctIF[321]  (.D(b4_nUAi[808]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[809]));
    SLE \b6_OKctIF[1064]  (.D(b4_nUAi[65]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[66]));
    SLE \b6_OKctIF[327]  (.D(b4_nUAi[802]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[803]));
    SLE \b6_OKctIF[133]  (.D(b4_nUAi[996]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[997]));
    SLE \b6_OKctIF[871]  (.D(b4_nUAi[258]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[259]));
    SLE \b6_OKctIF[603]  (.D(b4_nUAi[526]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[527]));
    SLE \b6_OKctIF[754]  (.D(b4_nUAi[375]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[376]));
    SLE \b6_OKctIF[735]  (.D(b4_nUAi[394]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[395]));
    SLE \b6_OKctIF[1109]  (.D(b4_nUAi[20]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[21]));
    SLE \b6_OKctIF[1117]  (.D(b4_nUAi[12]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[13]));
    SLE \b6_OKctIF[1079]  (.D(b4_nUAi[50]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[51]));
    SLE \b6_OKctIF[1008]  (.D(b4_nUAi[121]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[122]));
    SLE \b6_OKctIF[103]  (.D(b4_nUAi[1026]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1027]));
    SLE \b6_OKctIF[744]  (.D(b4_nUAi[385]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[386]));
    SLE \b6_OKctIF[156]  (.D(b4_nUAi[973]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[974]));
    SLE \b6_OKctIF[771]  (.D(b4_nUAi[358]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[359]));
    SLE \b6_OKctIF[705]  (.D(b4_nUAi[424]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[425]));
    VCC VCC (.Y(VCC_net_1));
    SLE \b6_OKctIF[923]  (.D(b4_nUAi[206]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[207]));
    SLE \b6_OKctIF[839]  (.D(b4_nUAi[290]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[291]));
    SLE \b6_OKctIF[146]  (.D(b4_nUAi[983]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[984]));
    SLE \b6_OKctIF[324]  (.D(b4_nUAi[805]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[806]));
    SLE \b6_OKctIF[517]  (.D(b4_nUAi[612]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[613]));
    SLE \b6_OKctIF[1010]  (.D(b4_nUAi[119]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[120]));
    SLE \b6_OKctIF[794]  (.D(b4_nUAi[335]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[336]));
    SLE \b6_OKctIF[114]  (.D(b4_nUAi[1015]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1016]));
    SLE \b6_OKctIF[939]  (.D(b4_nUAi[190]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[191]));
    SLE \b6_OKctIF[753]  (.D(b4_nUAi[376]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[377]));
    SLE \b6_OKctIF[562]  (.D(b4_nUAi[567]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[568]));
    SLE \b6_OKctIF[274]  (.D(b4_nUAi[855]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[856]));
    SLE \b6_OKctIF[809]  (.D(b4_nUAi[320]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[321]));
    SLE \b6_OKctIF[196]  (.D(b4_nUAi[933]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[934]));
    SLE \b6_OKctIF[858]  (.D(b4_nUAi[271]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[272]));
    SLE \b6_OKctIF[743]  (.D(b4_nUAi[386]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[387]));
    SLE \b6_OKctIF[253]  (.D(b4_nUAi[876]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[877]));
    SLE \b6_OKctIF[770]  (.D(b4_nUAi[359]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[360]));
    SLE \b6_OKctIF[581]  (.D(b4_nUAi[548]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[549]));
    SLE \b6_OKctIF[909]  (.D(b4_nUAi[220]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[221]));
    SLE \b6_OKctIF[1042]  (.D(b4_nUAi[87]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[88]));
    SLE \b6_OKctIF[937]  (.D(b4_nUAi[192]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[193]));
    SLE \b6_OKctIF[848]  (.D(b4_nUAi[281]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[282]));
    SLE \b6_OKctIF[243]  (.D(b4_nUAi[886]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[887]));
    SLE \b6_OKctIF[68]  (.D(b4_nUAi[1061]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1062]));
    SLE \b6_OKctIF[972]  (.D(b4_nUAi[157]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[158]));
    SLE \b6_OKctIF[834]  (.D(b4_nUAi[295]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[296]));
    SLE \b6_OKctIF[1046]  (.D(b4_nUAi[83]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[84]));
    SLE \b6_OKctIF[793]  (.D(b4_nUAi[336]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[337]));
    SLE \b6_OKctIF[729]  (.D(b4_nUAi[400]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[401]));
    SLE \b6_OKctIF[5]  (.D(b4_nUAi[1124]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1125]));
    SLE \b6_OKctIF[1055]  (.D(b4_nUAi[74]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[75]));
    SLE \b6_OKctIF[661]  (.D(b4_nUAi[468]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[469]));
    SLE \b6_OKctIF[555]  (.D(b4_nUAi[574]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[575]));
    SLE \b6_OKctIF[168]  (.D(b4_nUAi[961]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[962]));
    SLE \b6_OKctIF[438]  (.D(b4_nUAi[691]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[692]));
    SLE \b6_OKctIF[907]  (.D(b4_nUAi[222]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[223]));
    SLE \b6_OKctIF[489]  (.D(b4_nUAi[640]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[641]));
    SLE \b6_OKctIF[898]  (.D(b4_nUAi[231]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[232]));
    SLE \b6_OKctIF[293]  (.D(b4_nUAi[836]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[837]));
    SLE \b6_OKctIF[672]  (.D(b4_nUAi[457]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[458]));
    SLE \b6_OKctIF[867]  (.D(b4_nUAi[262]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[263]));
    SLE \b6_OKctIF[386]  (.D(b4_nUAi[743]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[744]));
    SLE \b6_OKctIF[804]  (.D(b4_nUAi[325]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[326]));
    SLE \b6_OKctIF[545]  (.D(b4_nUAi[584]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[585]));
    SLE \b6_OKctIF[637]  (.D(b4_nUAi[492]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[493]));
    SLE \b6_OKctIF[271]  (.D(b4_nUAi[858]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[859]));
    SLE \b6_OKctIF[408]  (.D(b4_nUAi[721]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[722]));
    SLE \b6_OKctIF[674]  (.D(b4_nUAi[455]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[456]));
    SLE \b6_OKctIF[466]  (.D(b4_nUAi[663]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[664]));
    SLE \b6_OKctIF[250]  (.D(b4_nUAi[879]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[880]));
    SLE \b6_OKctIF[956]  (.D(b4_nUAi[173]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[174]));
    SLE \b6_OKctIF[595]  (.D(b4_nUAi[534]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[535]));
    SLE \b6_OKctIF[318]  (.D(b4_nUAi[811]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[812]));
    SLE \b6_OKctIF[179]  (.D(b4_nUAi[950]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[951]));
    SLE \b6_OKctIF[607]  (.D(b4_nUAi[522]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[523]));
    SLE \b6_OKctIF[618]  (.D(b4_nUAi[511]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[512]));
    SLE \b6_OKctIF[823]  (.D(b4_nUAi[306]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[307]));
    SLE \b6_OKctIF[61]  (.D(b4_nUAi[1068]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1069]));
    SLE \b6_OKctIF[240]  (.D(b4_nUAi[889]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[890]));
    SLE \b6_OKctIF[946]  (.D(b4_nUAi[183]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[184]));
    SLE \b6_OKctIF[767]  (.D(b4_nUAi[362]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[363]));
    SLE \b6_OKctIF[911]  (.D(b4_nUAi[218]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[219]));
    SLE \b6_OKctIF[984]  (.D(b4_nUAi[145]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[146]));
    SLE \b6_OKctIF[856]  (.D(b4_nUAi[273]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[274]));
    SLE \b6_OKctIF[1108]  (.D(b4_nUAi[21]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[22]));
    SLE \b6_OKctIF[625]  (.D(b4_nUAi[504]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[505]));
    SLE \b6_OKctIF[18]  (.D(b4_nUAi[1111]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1112]));
    SLE \b6_OKctIF[55]  (.D(b4_nUAi[1074]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1075]));
    SLE \b6_OKctIF[290]  (.D(b4_nUAi[839]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[840]));
    SLE \b6_OKctIF[1061]  (.D(b4_nUAi[68]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[69]));
    SLE \b6_OKctIF[996]  (.D(b4_nUAi[133]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[134]));
    SLE \b6_OKctIF[50]  (.D(b4_nUAi[1079]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1080]));
    SLE \b6_OKctIF[846]  (.D(b4_nUAi[283]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[284]));
    SLE \b6_OKctIF[880]  (.D(b4_nUAi[249]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[250]));
    SLE \b6_OKctIF[120]  (.D(b4_nUAi[1009]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1010]));
    SLE \b6_OKctIF[1027]  (.D(b4_nUAi[102]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[103]));
    SLE \b6_OKctIF[568]  (.D(b4_nUAi[561]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[562]));
    SLE \b6_OKctIF[613]  (.D(b4_nUAi[516]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[517]));
    SLE \b6_OKctIF[451]  (.D(b4_nUAi[678]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[679]));
    SLE \b6_OKctIF[1023]  (.D(b4_nUAi[106]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[107]));
    SLE \b6_OKctIF[738]  (.D(b4_nUAi[391]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[392]));
    SLE \b6_OKctIF[896]  (.D(b4_nUAi[233]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[234]));
    SLE \b6_OKctIF[370]  (.D(b4_nUAi[759]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[760]));
    SLE \b6_OKctIF[113]  (.D(b4_nUAi[1016]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1017]));
    SLE \b6_OKctIF[1114]  (.D(b4_nUAi[15]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[16]));
    SLE \b6_OKctIF[361]  (.D(b4_nUAi[768]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[769]));
    SLE \b6_OKctIF[441]  (.D(b4_nUAi[688]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[689]));
    SLE \b6_OKctIF[367]  (.D(b4_nUAi[762]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[763]));
    SLE \b6_OKctIF[639]  (.D(b4_nUAi[490]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[491]));
    SLE \b6_OKctIF[98]  (.D(b4_nUAi[1031]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1032]));
    SLE \b6_OKctIF[715]  (.D(b4_nUAi[414]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[415]));
    SLE \b6_OKctIF[157]  (.D(b4_nUAi[972]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[973]));
    SLE \b6_OKctIF[1005]  (.D(b4_nUAi[124]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[125]));
    SLE \b6_OKctIF[708]  (.D(b4_nUAi[421]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[422]));
    SLE \b6_OKctIF[11]  (.D(b4_nUAi[1118]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1119]));
    SLE \b6_OKctIF[1069]  (.D(b4_nUAi[60]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[61]));
    SLE \b6_OKctIF[930]  (.D(b4_nUAi[199]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[200]));
    SLE \b6_OKctIF[491]  (.D(b4_nUAi[638]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[639]));
    SLE \b6_OKctIF[1110]  (.D(b4_nUAi[19]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[20]));
    SLE \b6_OKctIF[147]  (.D(b4_nUAi[982]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[983]));
    SLE \b6_OKctIF[609]  (.D(b4_nUAi[520]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[521]));
    SLE \b6_OKctIF[276]  (.D(b4_nUAi[853]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[854]));
    SLE \b6_OKctIF[520]  (.D(b4_nUAi[609]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[610]));
    SLE \b6_OKctIF[988]  (.D(b4_nUAi[141]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[142]));
    SLE \b6_OKctIF[228]  (.D(b4_nUAi[901]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[902]));
    SLE \b6_OKctIF[819]  (.D(b4_nUAi[310]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[311]));
    SLE \b6_OKctIF[474]  (.D(b4_nUAi[655]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[656]));
    SLE \b6_OKctIF[900]  (.D(b4_nUAi[229]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[230]));
    SLE \b6_OKctIF[963]  (.D(b4_nUAi[166]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[167]));
    SLE \b6_OKctIF[831]  (.D(b4_nUAi[298]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[299]));
    SLE \b6_OKctIF[197]  (.D(b4_nUAi[932]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[933]));
    SLE \b6_OKctIF[919]  (.D(b4_nUAi[210]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[211]));
    SLE \b6_OKctIF[584]  (.D(b4_nUAi[545]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[546]));
    SLE \b6_OKctIF[364]  (.D(b4_nUAi[765]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[766]));
    SLE \b6_OKctIF[91]  (.D(b4_nUAi[1038]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1039]));
    SLE \b6_OKctIF[589]  (.D(b4_nUAi[540]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[541]));
    SLE \b6_OKctIF[57]  (.D(b4_nUAi[1072]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1073]));
    SLE \b6_OKctIF[23]  (.D(b4_nUAi[1106]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1107]));
    SLE \b6_OKctIF[45]  (.D(b4_nUAi[1084]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1085]));
    SLE \b6_OKctIF[801]  (.D(b4_nUAi[328]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[329]));
    SLE \b6_OKctIF[40]  (.D(b4_nUAi[1089]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1090]));
    SLE \b6_OKctIF[917]  (.D(b4_nUAi[212]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[213]));
    SLE \b6_OKctIF[1084]  (.D(b4_nUAi[45]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[46]));
    SLE \b6_OKctIF[22]  (.D(b4_nUAi[1107]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1108]));
    SLE \b6_OKctIF[171]  (.D(b4_nUAi[958]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[959]));
    SLE \b6_OKctIF[814]  (.D(b4_nUAi[315]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[316]));
    SLE \b6_OKctIF[1127]  (.D(b4_nUAi[2]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[3]));
    SLE \b6_OKctIF[731]  (.D(b4_nUAi[398]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[399]));
    SLE \b6_OKctIF[54]  (.D(b4_nUAi[1075]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1076]));
    SLE \b6_OKctIF[523]  (.D(b4_nUAi[606]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[607]));
    SLE \b6_OKctIF[1101]  (.D(b4_nUAi[28]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[29]));
    SLE \b6_OKctIF[66]  (.D(b4_nUAi[1063]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1064]));
    SLE \b6_OKctIF[769]  (.D(b4_nUAi[360]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[361]));
    SLE \b6_OKctIF[418]  (.D(b4_nUAi[711]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[712]));
    SLE \b6_OKctIF[379]  (.D(b4_nUAi[750]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[751]));
    SLE \b6_OKctIF[422]  (.D(b4_nUAi[707]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[708]));
    SLE \b6_OKctIF[620]  (.D(b4_nUAi[509]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[510]));
    SLE \b6_OKctIF[59]  (.D(b4_nUAi[1070]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1071]));
    SLE \b6_OKctIF[701]  (.D(b4_nUAi[428]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[429]));
    SLE \b6_OKctIF[423]  (.D(b4_nUAi[706]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[707]));
    SLE \b6_OKctIF[0]  (.D(b4_nUAi[1129]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b7_PSyi3wy));
    SLE \b6_OKctIF[617]  (.D(b4_nUAi[512]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[513]));
    SLE \b6_OKctIF[234]  (.D(b4_nUAi[895]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[896]));
    SLE \b6_OKctIF[1020]  (.D(b4_nUAi[109]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[110]));
    SLE \b6_OKctIF[383]  (.D(b4_nUAi[746]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[747]));
    SLE \b6_OKctIF[730]  (.D(b4_nUAi[399]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[400]));
    SLE \b6_OKctIF[38]  (.D(b4_nUAi[1091]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1092]));
    SLE \b6_OKctIF[229]  (.D(b4_nUAi[900]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[901]));
    SLE \b6_OKctIF[287]  (.D(b4_nUAi[842]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[843]));
    SLE \b6_OKctIF[204]  (.D(b4_nUAi[925]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[926]));
    SLE \b6_OKctIF[932]  (.D(b4_nUAi[197]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[198]));
    SLE \b6_OKctIF[700]  (.D(b4_nUAi[429]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[430]));
    SLE \b6_OKctIF[73]  (.D(b4_nUAi[1056]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1057]));
    SLE \b6_OKctIF[863]  (.D(b4_nUAi[266]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[267]));
    SLE \b6_OKctIF[875]  (.D(b4_nUAi[254]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[255]));
    SLE \b6_OKctIF[632]  (.D(b4_nUAi[497]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[498]));
    SLE \b6_OKctIF[975]  (.D(b4_nUAi[154]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[155]));
    SLE \b6_OKctIF[72]  (.D(b4_nUAi[1057]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1058]));
    SLE \b6_OKctIF[902]  (.D(b4_nUAi[227]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[228]));
    SLE \b6_OKctIF[551]  (.D(b4_nUAi[578]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[579]));
    SLE \b6_OKctIF[665]  (.D(b4_nUAi[464]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[465]));
    SLE \b6_OKctIF[231]  (.D(b4_nUAi[898]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[899]));
    SLE \b6_OKctIF[16]  (.D(b4_nUAi[1113]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1114]));
    SLE \b6_OKctIF[634]  (.D(b4_nUAi[495]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[496]));
    SLE \b6_OKctIF[47]  (.D(b4_nUAi[1082]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1083]));
    SLE \b6_OKctIF[1038]  (.D(b4_nUAi[91]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[92]));
    SLE \b6_OKctIF[602]  (.D(b4_nUAi[527]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[528]));
    SLE \b6_OKctIF[541]  (.D(b4_nUAi[588]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[589]));
    SLE \b6_OKctIF[139]  (.D(b4_nUAi[990]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[991]));
    SLE \b6_OKctIF[31]  (.D(b4_nUAi[1098]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1099]));
    SLE \b6_OKctIF[160]  (.D(b4_nUAi[969]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[970]));
    SLE \b6_OKctIF[718]  (.D(b4_nUAi[411]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[412]));
    SLE \b6_OKctIF[44]  (.D(b4_nUAi[1085]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1086]));
    SLE \b6_OKctIF[459]  (.D(b4_nUAi[670]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[671]));
    SLE \b6_OKctIF[201]  (.D(b4_nUAi[928]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[929]));
    SLE \b6_OKctIF[604]  (.D(b4_nUAi[525]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[526]));
    SLE \b6_OKctIF[582]  (.D(b4_nUAi[547]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[548]));
    SLE \b6_OKctIF[356]  (.D(b4_nUAi[773]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[774]));
    SLE \b6_OKctIF[591]  (.D(b4_nUAi[538]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[539]));
    SLE \b6_OKctIF[122]  (.D(b4_nUAi[1007]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1008]));
    SLE \b6_OKctIF[619]  (.D(b4_nUAi[510]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[511]));
    SLE \b6_OKctIF[109]  (.D(b4_nUAi[1020]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1021]));
    SLE \b6_OKctIF[722]  (.D(b4_nUAi[407]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[408]));
    SLE \b6_OKctIF[449]  (.D(b4_nUAi[680]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[681]));
    SLE \b6_OKctIF[49]  (.D(b4_nUAi[1080]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1081]));
    SLE \b6_OKctIF[346]  (.D(b4_nUAi[783]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[784]));
    SLE \b6_OKctIF[275]  (.D(b4_nUAi[854]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[855]));
    SLE \b6_OKctIF[1113]  (.D(b4_nUAi[16]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[17]));
    SLE \b6_OKctIF[470]  (.D(b4_nUAi[659]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[660]));
    SLE \b6_OKctIF[96]  (.D(b4_nUAi[1033]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1034]));
    SLE \b6_OKctIF[1078]  (.D(b4_nUAi[51]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[52]));
    SLE \b6_OKctIF[372]  (.D(b4_nUAi[757]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[758]));
    SLE \b6_OKctIF[910]  (.D(b4_nUAi[219]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[220]));
    SLE \b6_OKctIF[1097]  (.D(b4_nUAi[32]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[33]));
    SLE \b6_OKctIF[499]  (.D(b4_nUAi[630]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[631]));
    SLE \b6_OKctIF[396]  (.D(b4_nUAi[733]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[734]));
    SLE \b6_OKctIF[1105]  (.D(b4_nUAi[24]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[25]));
    SLE \b6_OKctIF[1093]  (.D(b4_nUAi[36]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[37]));
    SLE \b6_OKctIF[560]  (.D(b4_nUAi[569]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[570]));
    SLE \b6_OKctIF[681]  (.D(b4_nUAi[448]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[449]));
    SLE \b6_OKctIF[188]  (.D(b4_nUAi[941]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[942]));
    SLE \b6_OKctIF[330]  (.D(b4_nUAi[799]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[800]));
    SLE \b6_OKctIF[268]  (.D(b4_nUAi[861]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[862]));
    SLE \b6_OKctIF[811]  (.D(b4_nUAi[318]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[319]));
    SLE \b6_OKctIF[1081]  (.D(b4_nUAi[48]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[49]));
    SLE \b6_OKctIF[887]  (.D(b4_nUAi[242]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[243]));
    SLE \b6_OKctIF[954]  (.D(b4_nUAi[175]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[176]));
    SLE \b6_OKctIF[1014]  (.D(b4_nUAi[115]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[116]));
    SLE \b6_OKctIF[425]  (.D(b4_nUAi[704]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[705]));
    SLE \b6_OKctIF[1124]  (.D(b4_nUAi[5]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[6]));
    SLE \b6_OKctIF[944]  (.D(b4_nUAi[185]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[186]));
    SLE \b6_OKctIF[822]  (.D(b4_nUAi[307]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[308]));
    SLE \b6_OKctIF[850]  (.D(b4_nUAi[279]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[280]));
    SLE \b6_OKctIF[300]  (.D(b4_nUAi[829]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[830]));
    SLE \b6_OKctIF[1112]  (.D(b4_nUAi[17]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[18]));
    SLE \b6_OKctIF[486]  (.D(b4_nUAi[643]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[644]));
    SLE \b6_OKctIF[9]  (.D(b4_nUAi[1120]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1121]));
    SLE \b6_OKctIF[626]  (.D(b4_nUAi[503]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[504]));
    SLE \b6_OKctIF[236]  (.D(b4_nUAi[893]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[894]));
    SLE \b6_OKctIF[840]  (.D(b4_nUAi[289]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[290]));
    SLE \b6_OKctIF[726]  (.D(b4_nUAi[403]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[404]));
    SLE \b6_OKctIF[711]  (.D(b4_nUAi[418]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[419]));
    SLE \b6_OKctIF[994]  (.D(b4_nUAi[135]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[136]));
    SLE \b6_OKctIF[427]  (.D(b4_nUAi[702]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[703]));
    SLE \b6_OKctIF[1106]  (.D(b4_nUAi[23]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[24]));
    SLE \b6_OKctIF[1120]  (.D(b4_nUAi[9]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[10]));
    SLE \b6_OKctIF[434]  (.D(b4_nUAi[695]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[696]));
    SLE \b6_OKctIF[787]  (.D(b4_nUAi[342]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[343]));
    SLE \b6_OKctIF[563]  (.D(b4_nUAi[566]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[567]));
    SLE \b6_OKctIF[1052]  (.D(b4_nUAi[77]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[78]));
    SLE \b6_OKctIF[890]  (.D(b4_nUAi[239]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[240]));
    SLE \b6_OKctIF[206]  (.D(b4_nUAi[923]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[924]));
    SLE \b6_OKctIF[1089]  (.D(b4_nUAi[40]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[41]));
    SLE \b6_OKctIF[325]  (.D(b4_nUAi[804]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[805]));
    SLE \b6_OKctIF[462]  (.D(b4_nUAi[667]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[668]));
    SLE \b6_OKctIF[214]  (.D(b4_nUAi[915]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[916]));
    SLE \b6_OKctIF[660]  (.D(b4_nUAi[469]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[470]));
    SLE \b6_OKctIF[1056]  (.D(b4_nUAi[73]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[74]));
    SLE \b6_OKctIF[774]  (.D(b4_nUAi[355]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[356]));
    SLE \b6_OKctIF[404]  (.D(b4_nUAi[725]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[726]));
    SLE \b6_OKctIF[710]  (.D(b4_nUAi[419]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[420]));
    SLE \b6_OKctIF[463]  (.D(b4_nUAi[666]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[667]));
    SLE \b6_OKctIF[588]  (.D(b4_nUAi[541]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[542]));
    SLE \b6_OKctIF[958]  (.D(b4_nUAi[171]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[172]));
    SLE \b6_OKctIF[176]  (.D(b4_nUAi[953]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[954]));
    SLE \b6_OKctIF[131]  (.D(b4_nUAi[998]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[999]));
    SLE \b6_OKctIF[912]  (.D(b4_nUAi[217]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[218]));
    SLE \b6_OKctIF[36]  (.D(b4_nUAi[1093]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1094]));
    SLE \b6_OKctIF[222]  (.D(b4_nUAi[907]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[908]));
    SLE \b6_OKctIF[948]  (.D(b4_nUAi[181]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[182]));
    SLE \b6_OKctIF[269]  (.D(b4_nUAi[860]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[861]));
    SLE \b6_OKctIF[554]  (.D(b4_nUAi[575]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[576]));
    SLE \b6_OKctIF[381]  (.D(b4_nUAi[748]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[749]));
    SLE \b6_OKctIF[387]  (.D(b4_nUAi[742]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[743]));
    SLE \b6_OKctIF[339]  (.D(b4_nUAi[790]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[791]));
    SLE \b6_OKctIF[125]  (.D(b4_nUAi[1004]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1005]));
    SLE \b6_OKctIF[526]  (.D(b4_nUAi[603]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[604]));
    SLE \b6_OKctIF[612]  (.D(b4_nUAi[517]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[518]));
    SLE \b6_OKctIF[101]  (.D(b4_nUAi[1028]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1029]));
    SLE \b6_OKctIF[773]  (.D(b4_nUAi[356]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[357]));
    SLE \b6_OKctIF[544]  (.D(b4_nUAi[585]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[586]));
    SLE \b6_OKctIF[559]  (.D(b4_nUAi[570]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[571]));
    SLE \b6_OKctIF[1090]  (.D(b4_nUAi[39]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[40]));
    SLE \b6_OKctIF[998]  (.D(b4_nUAi[131]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[132]));
    SLE \b6_OKctIF[878]  (.D(b4_nUAi[251]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[252]));
    SLE \b6_OKctIF[273]  (.D(b4_nUAi[856]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[857]));
    SLE \b6_OKctIF[211]  (.D(b4_nUAi[918]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[919]));
    SLE \b6_OKctIF[1035]  (.D(b4_nUAi[94]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[95]));
    SLE \b6_OKctIF[309]  (.D(b4_nUAi[820]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[821]));
    SLE \b6_OKctIF[614]  (.D(b4_nUAi[515]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[516]));
    SLE \b6_OKctIF[549]  (.D(b4_nUAi[580]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[581]));
    SLE \b6_OKctIF[594]  (.D(b4_nUAi[535]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[536]));
    SLE \b6_OKctIF[119]  (.D(b4_nUAi[1010]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1011]));
    SLE \b6_OKctIF[983]  (.D(b4_nUAi[146]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[147]));
    SLE \b6_OKctIF[599]  (.D(b4_nUAi[530]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[531]));
    SLE \b6_OKctIF[25]  (.D(b4_nUAi[1104]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1105]));
    SLE \b6_OKctIF[384]  (.D(b4_nUAi[745]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[746]));
    SLE \b6_OKctIF[575]  (.D(b4_nUAi[554]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[555]));
    SLE \b6_OKctIF[20]  (.D(b4_nUAi[1109]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1110]));
    SLE \b6_OKctIF[835]  (.D(b4_nUAi[294]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[295]));
    SLE \b6_OKctIF[935]  (.D(b4_nUAi[194]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[195]));
    SLE \b6_OKctIF[527]  (.D(b4_nUAi[602]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[603]));
    SLE \b6_OKctIF[353]  (.D(b4_nUAi[776]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[777]));
    SLE \b6_OKctIF[162]  (.D(b4_nUAi[967]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[968]));
    SLE \b6_OKctIF[124]  (.D(b4_nUAi[1005]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1006]));
    SLE \b6_OKctIF[1075]  (.D(b4_nUAi[54]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[55]));
    SLE \b6_OKctIF[762]  (.D(b4_nUAi[367]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[368]));
    SLE \b6_OKctIF[1068]  (.D(b4_nUAi[61]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[62]));
    SLE \b6_OKctIF[1002]  (.D(b4_nUAi[127]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[128]));
    SLE \b6_OKctIF[805]  (.D(b4_nUAi[324]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[325]));
    SLE \b6_OKctIF[343]  (.D(b4_nUAi[786]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[787]));
    SLE \b6_OKctIF[1011]  (.D(b4_nUAi[118]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[119]));
    SLE \b6_OKctIF[257]  (.D(b4_nUAi[872]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[873]));
    SLE \b6_OKctIF[270]  (.D(b4_nUAi[859]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[860]));
    SLE \b6_OKctIF[905]  (.D(b4_nUAi[224]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[225]));
    SLE \b6_OKctIF[1006]  (.D(b4_nUAi[123]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[124]));
    SLE \b6_OKctIF[976]  (.D(b4_nUAi[153]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[154]));
    
endmodule


module b8_1LbcQDr1_x_85_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [291:291] mdiclink_reg;
input  [85:85] b11_OFWNT9L_8tZ;
input  [875:873] b4_nUAi;
output [291:291] b6_2ZTGIf;

    wire b3_P_F_6_bm_105, b3_P_F_6_am_105, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_105), .B(
        b4_nUAi[875]), .C(b3_P_F_6_am_105), .Y(b6_2ZTGIf[291]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[291]), .B(
        b11_OFWNT9L_8tZ[85]), .C(b4_nUAi[874]), .D(b4_nUAi[873]), .Y(
        b3_P_F_6_am_105));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[291]), .B(
        b11_OFWNT9L_8tZ[85]), .C(b4_nUAi[873]), .D(b4_nUAi[874]), .Y(
        b3_P_F_6_bm_105));
    
endmodule


module b8_1LbcQDr1_x_69_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [307:307] mdiclink_reg;
input  [69:69] b11_OFWNT9L_8tZ;
input  [923:921] b4_nUAi;
output [307:307] b6_2ZTGIf;

    wire b3_P_F_6_bm_115, b3_P_F_6_am_115, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_115), .B(
        b4_nUAi[923]), .C(b3_P_F_6_am_115), .Y(b6_2ZTGIf[307]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[307]), .B(
        b11_OFWNT9L_8tZ[69]), .C(b4_nUAi[922]), .D(b4_nUAi[921]), .Y(
        b3_P_F_6_am_115));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[307]), .B(
        b11_OFWNT9L_8tZ[69]), .C(b4_nUAi[921]), .D(b4_nUAi[922]), .Y(
        b3_P_F_6_bm_115));
    
endmodule


module b8_1LbcQDr1_x_16_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [360:360] mdiclink_reg;
input  [16:16] b11_OFWNT9L_8tZ;
input  [1082:1080] b4_nUAi;
output [360:360] b6_2ZTGIf;

    wire b3_P_F_6_bm_141, b3_P_F_6_am_141, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_141), .B(
        b4_nUAi[1082]), .C(b3_P_F_6_am_141), .Y(b6_2ZTGIf[360]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[360]), .B(
        b11_OFWNT9L_8tZ[16]), .C(b4_nUAi[1081]), .D(b4_nUAi[1080]), .Y(
        b3_P_F_6_am_141));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[360]), .B(
        b11_OFWNT9L_8tZ[16]), .C(b4_nUAi[1080]), .D(b4_nUAi[1081]), .Y(
        b3_P_F_6_bm_141));
    
endmodule


module b8_1LbcQDr1_x_248_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [128:128] mdiclink_reg;
input  [248:248] b11_OFWNT9L_8tZ;
input  [386:384] b4_nUAi;
output [128:128] b6_2ZTGIf;

    wire b3_P_F_6_bm_28, b3_P_F_6_am_28, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_28), .B(
        b4_nUAi[386]), .C(b3_P_F_6_am_28), .Y(b6_2ZTGIf[128]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[128]), .B(
        b11_OFWNT9L_8tZ[248]), .C(b4_nUAi[385]), .D(b4_nUAi[384]), .Y(
        b3_P_F_6_am_28));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[128]), .B(
        b11_OFWNT9L_8tZ[248]), .C(b4_nUAi[384]), .D(b4_nUAi[385]), .Y(
        b3_P_F_6_bm_28));
    
endmodule


module b8_1LbcQDr1_x_32_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [344:344] mdiclink_reg;
input  [32:32] b11_OFWNT9L_8tZ;
input  [1034:1032] b4_nUAi;
output [344:344] b6_2ZTGIf;

    wire b3_P_F_6_bm_131, b3_P_F_6_am_131, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_131), .B(
        b4_nUAi[1034]), .C(b3_P_F_6_am_131), .Y(b6_2ZTGIf[344]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[344]), .B(
        b11_OFWNT9L_8tZ[32]), .C(b4_nUAi[1033]), .D(b4_nUAi[1032]), .Y(
        b3_P_F_6_am_131));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[344]), .B(
        b11_OFWNT9L_8tZ[32]), .C(b4_nUAi[1032]), .D(b4_nUAi[1033]), .Y(
        b3_P_F_6_bm_131));
    
endmodule


module b8_1LbcQDr1_x_302_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [74:74] mdiclink_reg;
input  [302:302] b11_OFWNT9L_8tZ;
input  [224:222] b4_nUAi;
output [74:74] b6_2ZTGIf;

    wire b3_P_F_6_bm_193, b3_P_F_6_am_193, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_193), .B(
        b4_nUAi[224]), .C(b3_P_F_6_am_193), .Y(b6_2ZTGIf[74]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[74]), .B(
        b11_OFWNT9L_8tZ[302]), .C(b4_nUAi[223]), .D(b4_nUAi[222]), .Y(
        b3_P_F_6_am_193));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[74]), .B(
        b11_OFWNT9L_8tZ[302]), .C(b4_nUAi[222]), .D(b4_nUAi[223]), .Y(
        b3_P_F_6_bm_193));
    
endmodule


module b8_1LbcQDr1_x_136_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [240:240] mdiclink_reg;
input  [136:136] b11_OFWNT9L_8tZ;
input  [722:720] b4_nUAi;
output [240:240] b6_2ZTGIf;

    wire b3_P_F_6_bm_232, b3_P_F_6_am_232, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_232), .B(
        b4_nUAi[722]), .C(b3_P_F_6_am_232), .Y(b6_2ZTGIf[240]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[240]), .B(
        b11_OFWNT9L_8tZ[136]), .C(b4_nUAi[721]), .D(b4_nUAi[720]), .Y(
        b3_P_F_6_am_232));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[240]), .B(
        b11_OFWNT9L_8tZ[136]), .C(b4_nUAi[720]), .D(b4_nUAi[721]), .Y(
        b3_P_F_6_bm_232));
    
endmodule


module b8_1LbcQDr1_x_225_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [151:151] mdiclink_reg;
input  [225:225] b11_OFWNT9L_8tZ;
input  [455:453] b4_nUAi;
output [151:151] b6_2ZTGIf;

    wire b3_P_F_6_bm_32, b3_P_F_6_am_32, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_32), .B(
        b4_nUAi[455]), .C(b3_P_F_6_am_32), .Y(b6_2ZTGIf[151]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[151]), .B(
        b11_OFWNT9L_8tZ[225]), .C(b4_nUAi[454]), .D(b4_nUAi[453]), .Y(
        b3_P_F_6_am_32));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[151]), .B(
        b11_OFWNT9L_8tZ[225]), .C(b4_nUAi[453]), .D(b4_nUAi[454]), .Y(
        b3_P_F_6_bm_32));
    
endmodule


module b8_1LbcQDr1_x_183_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [193:193] mdiclink_reg;
input  [183:183] b11_OFWNT9L_8tZ;
input  [581:579] b4_nUAi;
output [193:193] b6_2ZTGIf;

    wire b3_P_F_6_bm_67, b3_P_F_6_am_67, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_67), .B(
        b4_nUAi[581]), .C(b3_P_F_6_am_67), .Y(b6_2ZTGIf[193]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[193]), .B(
        b11_OFWNT9L_8tZ[183]), .C(b4_nUAi[580]), .D(b4_nUAi[579]), .Y(
        b3_P_F_6_am_67));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[193]), .B(
        b11_OFWNT9L_8tZ[183]), .C(b4_nUAi[579]), .D(b4_nUAi[580]), .Y(
        b3_P_F_6_bm_67));
    
endmodule


module b8_1LbcQDr1_x_249_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [127:127] mdiclink_reg;
input  [249:249] b11_OFWNT9L_8tZ;
input  [382:381] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[127]), .B(
        b11_OFWNT9L_8tZ[249]), .C(b4_nUAi[382]), .D(b4_nUAi[381]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[127]), .B(
        b11_OFWNT9L_8tZ[249]), .C(b4_nUAi[382]), .D(b4_nUAi[381]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_362_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [14:14] mdiclink_reg;
input  [362:362] b11_OFWNT9L_8tZ;
input  [43:42] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[14]), .B(
        b11_OFWNT9L_8tZ[362]), .C(b4_nUAi[43]), .D(b4_nUAi[42]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[14]), .B(
        b11_OFWNT9L_8tZ[362]), .C(b4_nUAi[43]), .D(b4_nUAi[42]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_164_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [212:212] mdiclink_reg;
input  [164:164] b11_OFWNT9L_8tZ;
input  [638:636] b4_nUAi;
output [212:212] b6_2ZTGIf;

    wire b3_P_F_6_bm_74, b3_P_F_6_am_74, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_74), .B(
        b4_nUAi[638]), .C(b3_P_F_6_am_74), .Y(b6_2ZTGIf[212]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[212]), .B(
        b11_OFWNT9L_8tZ[164]), .C(b4_nUAi[637]), .D(b4_nUAi[636]), .Y(
        b3_P_F_6_am_74));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[212]), .B(
        b11_OFWNT9L_8tZ[164]), .C(b4_nUAi[636]), .D(b4_nUAi[637]), .Y(
        b3_P_F_6_bm_74));
    
endmodule


module b8_1LbcQDr1_x_143_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [233:233] mdiclink_reg;
input  [143:143] b11_OFWNT9L_8tZ;
input  [701:699] b4_nUAi;
output [233:233] b6_2ZTGIf;

    wire b3_P_F_6_bm_214, b3_P_F_6_am_214, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_214), .B(
        b4_nUAi[701]), .C(b3_P_F_6_am_214), .Y(b6_2ZTGIf[233]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[233]), .B(
        b11_OFWNT9L_8tZ[143]), .C(b4_nUAi[700]), .D(b4_nUAi[699]), .Y(
        b3_P_F_6_am_214));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[233]), .B(
        b11_OFWNT9L_8tZ[143]), .C(b4_nUAi[699]), .D(b4_nUAi[700]), .Y(
        b3_P_F_6_bm_214));
    
endmodule


module b8_1LbcQDr1_x_36_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [340:340] mdiclink_reg;
input  [36:36] b11_OFWNT9L_8tZ;
input  [1022:1020] b4_nUAi;
output [340:340] b6_2ZTGIf;

    wire b3_P_F_6_bm_134, b3_P_F_6_am_134, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_134), .B(
        b4_nUAi[1022]), .C(b3_P_F_6_am_134), .Y(b6_2ZTGIf[340]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[340]), .B(
        b11_OFWNT9L_8tZ[36]), .C(b4_nUAi[1021]), .D(b4_nUAi[1020]), .Y(
        b3_P_F_6_am_134));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[340]), .B(
        b11_OFWNT9L_8tZ[36]), .C(b4_nUAi[1020]), .D(b4_nUAi[1021]), .Y(
        b3_P_F_6_bm_134));
    
endmodule


module b8_1LbcQDr1_x_24_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [352:352] mdiclink_reg;
input  [24:24] b11_OFWNT9L_8tZ;
input  [1058:1056] b4_nUAi;
output [352:352] b6_2ZTGIf;

    wire b3_P_F_6_bm_148, b3_P_F_6_am_148, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_148), .B(
        b4_nUAi[1058]), .C(b3_P_F_6_am_148), .Y(b6_2ZTGIf[352]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[352]), .B(
        b11_OFWNT9L_8tZ[24]), .C(b4_nUAi[1057]), .D(b4_nUAi[1056]), .Y(
        b3_P_F_6_am_148));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[352]), .B(
        b11_OFWNT9L_8tZ[24]), .C(b4_nUAi[1056]), .D(b4_nUAi[1057]), .Y(
        b3_P_F_6_bm_148));
    
endmodule


module b8_1LbcQDr1_x_174_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [202:202] mdiclink_reg;
input  [174:174] b11_OFWNT9L_8tZ;
input  [608:606] b4_nUAi;
output [202:202] b6_2ZTGIf;

    wire b3_P_F_6_bm_59, b3_P_F_6_am_59, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_59), .B(
        b4_nUAi[608]), .C(b3_P_F_6_am_59), .Y(b6_2ZTGIf[202]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[202]), .B(
        b11_OFWNT9L_8tZ[174]), .C(b4_nUAi[607]), .D(b4_nUAi[606]), .Y(
        b3_P_F_6_am_59));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[202]), .B(
        b11_OFWNT9L_8tZ[174]), .C(b4_nUAi[606]), .D(b4_nUAi[607]), .Y(
        b3_P_F_6_bm_59));
    
endmodule


module b8_1LbcQDr1_x_305_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [71:71] mdiclink_reg;
input  [305:305] b11_OFWNT9L_8tZ;
input  [215:213] b4_nUAi;
output [71:71] b6_2ZTGIf;

    wire b3_P_F_6_bm_196, b3_P_F_6_am_196, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_196), .B(
        b4_nUAi[215]), .C(b3_P_F_6_am_196), .Y(b6_2ZTGIf[71]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[71]), .B(
        b11_OFWNT9L_8tZ[305]), .C(b4_nUAi[214]), .D(b4_nUAi[213]), .Y(
        b3_P_F_6_am_196));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[71]), .B(
        b11_OFWNT9L_8tZ[305]), .C(b4_nUAi[213]), .D(b4_nUAi[214]), .Y(
        b3_P_F_6_bm_196));
    
endmodule


module b8_1LbcQDr1_x_365_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [11:11] mdiclink_reg;
input  [365:365] b11_OFWNT9L_8tZ;
input  [34:33] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[11]), .B(
        b11_OFWNT9L_8tZ[365]), .C(b4_nUAi[34]), .D(b4_nUAi[33]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[11]), .B(
        b11_OFWNT9L_8tZ[365]), .C(b4_nUAi[34]), .D(b4_nUAi[33]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_256_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [120:120] mdiclink_reg;
input  [256:256] b11_OFWNT9L_8tZ;
input  [362:360] b4_nUAi;
output [120:120] b6_2ZTGIf;

    wire b3_P_F_6_bm_11, b3_P_F_6_am_11, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_11), .B(
        b4_nUAi[362]), .C(b3_P_F_6_am_11), .Y(b6_2ZTGIf[120]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[120]), .B(
        b11_OFWNT9L_8tZ[256]), .C(b4_nUAi[361]), .D(b4_nUAi[360]), .Y(
        b3_P_F_6_am_11));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[120]), .B(
        b11_OFWNT9L_8tZ[256]), .C(b4_nUAi[360]), .D(b4_nUAi[361]), .Y(
        b3_P_F_6_bm_11));
    
endmodule


module b8_1LbcQDr1_x_101_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [275:275] mdiclink_reg;
input  [101:101] b11_OFWNT9L_8tZ;
input  [827:825] b4_nUAi;
output [275:275] b6_2ZTGIf;

    wire b3_P_F_6_bm_95, b3_P_F_6_am_95, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_95), .B(
        b4_nUAi[827]), .C(b3_P_F_6_am_95), .Y(b6_2ZTGIf[275]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[275]), .B(
        b11_OFWNT9L_8tZ[101]), .C(b4_nUAi[826]), .D(b4_nUAi[825]), .Y(
        b3_P_F_6_am_95));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[275]), .B(
        b11_OFWNT9L_8tZ[101]), .C(b4_nUAi[825]), .D(b4_nUAi[826]), .Y(
        b3_P_F_6_bm_95));
    
endmodule


module b8_1LbcQDr1_x_306_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [70:70] mdiclink_reg;
input  [306:306] b11_OFWNT9L_8tZ;
input  [212:210] b4_nUAi;
output [70:70] b6_2ZTGIf;

    wire b3_P_F_6_bm_197, b3_P_F_6_am_197, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_197), .B(
        b4_nUAi[212]), .C(b3_P_F_6_am_197), .Y(b6_2ZTGIf[70]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[70]), .B(
        b11_OFWNT9L_8tZ[306]), .C(b4_nUAi[211]), .D(b4_nUAi[210]), .Y(
        b3_P_F_6_am_197));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[70]), .B(
        b11_OFWNT9L_8tZ[306]), .C(b4_nUAi[210]), .D(b4_nUAi[211]), .Y(
        b3_P_F_6_bm_197));
    
endmodule


module b8_1LbcQDr1_x_366_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [10:10] mdiclink_reg;
input  [366:366] b11_OFWNT9L_8tZ;
input  [32:30] b4_nUAi;
output [10:10] b6_2ZTGIf;

    wire b3_P_F_6_bm_153, b3_P_F_6_am_153, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_153), .B(
        b4_nUAi[32]), .C(b3_P_F_6_am_153), .Y(b6_2ZTGIf[10]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[10]), .B(
        b11_OFWNT9L_8tZ[366]), .C(b4_nUAi[31]), .D(b4_nUAi[30]), .Y(
        b3_P_F_6_am_153));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[10]), .B(
        b11_OFWNT9L_8tZ[366]), .C(b4_nUAi[30]), .D(b4_nUAi[31]), .Y(
        b3_P_F_6_bm_153));
    
endmodule


module b8_1LbcQDr1_x_204_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [172:172] mdiclink_reg;
input  [204:204] b11_OFWNT9L_8tZ;
input  [517:516] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[172]), .B(
        b11_OFWNT9L_8tZ[204]), .C(b4_nUAi[517]), .D(b4_nUAi[516]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[172]), .B(
        b11_OFWNT9L_8tZ[204]), .C(b4_nUAi[517]), .D(b4_nUAi[516]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_325_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [51:51] mdiclink_reg;
input  [325:325] b11_OFWNT9L_8tZ;
input  [155:153] b4_nUAi;
output [51:51] b6_2ZTGIf;

    wire b3_P_F_6_bm_189, b3_P_F_6_am_189, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_189), .B(
        b4_nUAi[155]), .C(b3_P_F_6_am_189), .Y(b6_2ZTGIf[51]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[51]), .B(
        b11_OFWNT9L_8tZ[325]), .C(b4_nUAi[154]), .D(b4_nUAi[153]), .Y(
        b3_P_F_6_am_189));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[51]), .B(
        b11_OFWNT9L_8tZ[325]), .C(b4_nUAi[153]), .D(b4_nUAi[154]), .Y(
        b3_P_F_6_bm_189));
    
endmodule


module b9_O2yyf_fG2_x_22_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [10:10] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[10]));
    
endmodule


module b9_O2yyf_fG2_x_17_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [15:15] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[15]));
    
endmodule


module b9_O2yyf_fG2_x_14_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [18:18] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[18]));
    
endmodule


module b9_O2yyf_fG2_x_29_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [3:3] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[3]));
    
endmodule


module b9_O2yyf_fG2_x_19_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [13:13] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[13]));
    
endmodule


module b9_O2yyf_fG2_x_26_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [6:6] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[6]));
    
endmodule


module b9_O2yyf_fG2_x_12_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [20:20] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[20]));
    
endmodule


module b9_O2yyf_fG2_x_9_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_18,
       b4_nUAi_12,
       b4_nUAi_6,
       b4_nUAi_0,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_2,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       b7_PSyi3wy,
       N_27_3
    );
output [23:23] b13_CZS0wfY_d_FH9;
input  b4_nUAi_18;
input  b4_nUAi_12;
input  b4_nUAi_6;
input  b4_nUAi_0;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  b7_PSyi3wy;
input  N_27_3;

    wire o_3_net_1, o_2_net_1, o_1_net_1, o_0_net_1, o_4_net_1, 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_0), .B(b4_nUAi_12), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_1), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_2), .D(N_27_1), .Y(o_1_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_3), .B(b7_PSyi3wy), .C(
        o_0_net_1), .D(N_27_3), .Y(o_4_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_3_net_1));
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_2), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_0), .D(N_27_2), .Y(o_0_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_1_net_1), .B(o_4_net_1), .C(
        o_3_net_1), .D(o_2_net_1), .Y(b13_CZS0wfY_d_FH9[23]));
    GND GND (.Y(GND_net_1));
    
endmodule


module b9_O2yyf_fG2_x_16_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [16:16] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[16]));
    
endmodule


module b9_O2yyf_fG2_x_20_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [12:12] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[12]));
    
endmodule


module b9_O2yyf_fG2_x_21_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [11:11] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[11]));
    
endmodule


module b9_O2yyf_fG2_x_32_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [0:0] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[0]));
    
endmodule


module b9_O2yyf_fG2_x_31_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [1:1] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[1]));
    
endmodule


module b9_O2yyf_fG2_x_0_0(
       b14_CZS0wfY_d_FH9m,
       b11_uUT0JC4gFrY
    );
input  [23:0] b14_CZS0wfY_d_FH9m;
output [1:1] b11_uUT0JC4gFrY;

    wire o_17_net_1, o_16_net_1, o_15_net_1, o_14_net_1, o_13_net_1, 
        o_12_net_1, o_21_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h8000) )  o_16 (.A(b14_CZS0wfY_d_FH9m[11]), .B(
        b14_CZS0wfY_d_FH9m[10]), .C(b14_CZS0wfY_d_FH9m[9]), .D(
        b14_CZS0wfY_d_FH9m[8]), .Y(o_16_net_1));
    CFG4 #( .INIT(16'h8000) )  o_14 (.A(b14_CZS0wfY_d_FH9m[3]), .B(
        b14_CZS0wfY_d_FH9m[2]), .C(b14_CZS0wfY_d_FH9m[1]), .D(
        b14_CZS0wfY_d_FH9m[0]), .Y(o_14_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(b14_CZS0wfY_d_FH9m[19]), .B(
        b14_CZS0wfY_d_FH9m[18]), .C(b14_CZS0wfY_d_FH9m[17]), .D(
        b14_CZS0wfY_d_FH9m[16]), .Y(o_12_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h80) )  o (.A(o_16_net_1), .B(o_21_net_1), .C(
        o_17_net_1), .Y(b11_uUT0JC4gFrY[1]));
    CFG4 #( .INIT(16'h8000) )  o_17 (.A(b14_CZS0wfY_d_FH9m[15]), .B(
        b14_CZS0wfY_d_FH9m[14]), .C(b14_CZS0wfY_d_FH9m[13]), .D(
        b14_CZS0wfY_d_FH9m[12]), .Y(o_17_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h8000) )  o_13 (.A(b14_CZS0wfY_d_FH9m[23]), .B(
        b14_CZS0wfY_d_FH9m[22]), .C(b14_CZS0wfY_d_FH9m[21]), .D(
        b14_CZS0wfY_d_FH9m[20]), .Y(o_13_net_1));
    CFG4 #( .INIT(16'h8000) )  o_21 (.A(o_15_net_1), .B(o_14_net_1), 
        .C(o_13_net_1), .D(o_12_net_1), .Y(o_21_net_1));
    CFG4 #( .INIT(16'h8000) )  o_15 (.A(b14_CZS0wfY_d_FH9m[7]), .B(
        b14_CZS0wfY_d_FH9m[6]), .C(b14_CZS0wfY_d_FH9m[5]), .D(
        b14_CZS0wfY_d_FH9m[4]), .Y(o_15_net_1));
    
endmodule


module b9_O2yyf_fG2_x_27_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [5:5] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[5]));
    
endmodule


module b9_O2yyf_fG2_x_28_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [4:4] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[4]));
    
endmodule


module b9_O2yyf_fG2_x_10_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [22:22] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[22]));
    
endmodule


module b9_O2yyf_fG2_x_11_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [21:21] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[21]));
    
endmodule


module b9_O2yyf_fG2_x_24_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [8:8] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[8]));
    
endmodule


module b9_O2yyf_fG2_x_13_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [19:19] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[19]));
    
endmodule


module b9_O2yyf_fG2_x_15_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [17:17] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[17]));
    
endmodule


module b9_O2yyf_fG2_x_18_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [14:14] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[14]));
    
endmodule


module b9_O2yyf_fG2_x_30_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [2:2] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[2]));
    
endmodule


module b9_O2yyf_fG2_x_25_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [7:7] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[7]));
    
endmodule


module b9_O2yyf_fG2_x_23_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [9:9] b13_CZS0wfY_d_FH9;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_18), .C(
        b6_2ZTGIf_0), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_27), .C(
        b6_2ZTGIf_3), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_7), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_21), .C(
        b6_2ZTGIf_1), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_2), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_6), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_4), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[9]));
    
endmodule


module b16_CRGcTCua_eH4_2j7_x_0(
       b11_uUT0JC4gFrY,
       b4_nUAi_0,
       b4_nUAi_30,
       b4_nUAi_27,
       b4_nUAi_24,
       b4_nUAi_21,
       b4_nUAi_18,
       b4_nUAi_48,
       b4_nUAi_78,
       b4_nUAi_75,
       b4_nUAi_72,
       b4_nUAi_69,
       b4_nUAi_66,
       b4_nUAi_96,
       b4_nUAi_126,
       b4_nUAi_123,
       b4_nUAi_120,
       b4_nUAi_117,
       b4_nUAi_114,
       b4_nUAi_144,
       b4_nUAi_174,
       b4_nUAi_171,
       b4_nUAi_168,
       b4_nUAi_165,
       b4_nUAi_162,
       b4_nUAi_192,
       b4_nUAi_222,
       b4_nUAi_219,
       b4_nUAi_216,
       b4_nUAi_213,
       b4_nUAi_210,
       b4_nUAi_240,
       b4_nUAi_270,
       b4_nUAi_267,
       b4_nUAi_264,
       b4_nUAi_261,
       b4_nUAi_258,
       b4_nUAi_288,
       b4_nUAi_318,
       b4_nUAi_315,
       b4_nUAi_312,
       b4_nUAi_309,
       b4_nUAi_306,
       b4_nUAi_336,
       b4_nUAi_366,
       b4_nUAi_363,
       b4_nUAi_360,
       b4_nUAi_357,
       b4_nUAi_354,
       b4_nUAi_384,
       b4_nUAi_414,
       b4_nUAi_411,
       b4_nUAi_408,
       b4_nUAi_405,
       b4_nUAi_402,
       b4_nUAi_432,
       b4_nUAi_462,
       b4_nUAi_459,
       b4_nUAi_456,
       b4_nUAi_453,
       b4_nUAi_450,
       b4_nUAi_480,
       b4_nUAi_510,
       b4_nUAi_507,
       b4_nUAi_504,
       b4_nUAi_501,
       b4_nUAi_498,
       b4_nUAi_528,
       b4_nUAi_558,
       b4_nUAi_555,
       b4_nUAi_552,
       b4_nUAi_549,
       b4_nUAi_546,
       b4_nUAi_576,
       b4_nUAi_606,
       b4_nUAi_603,
       b4_nUAi_600,
       b4_nUAi_597,
       b4_nUAi_594,
       b4_nUAi_624,
       b4_nUAi_654,
       b4_nUAi_651,
       b4_nUAi_648,
       b4_nUAi_645,
       b4_nUAi_642,
       b4_nUAi_672,
       b4_nUAi_702,
       b4_nUAi_699,
       b4_nUAi_696,
       b4_nUAi_693,
       b4_nUAi_690,
       b4_nUAi_720,
       b4_nUAi_750,
       b4_nUAi_747,
       b4_nUAi_744,
       b4_nUAi_741,
       b4_nUAi_738,
       b4_nUAi_768,
       b4_nUAi_798,
       b4_nUAi_795,
       b4_nUAi_792,
       b4_nUAi_789,
       b4_nUAi_786,
       b4_nUAi_816,
       b4_nUAi_846,
       b4_nUAi_843,
       b4_nUAi_840,
       b4_nUAi_837,
       b4_nUAi_834,
       b4_nUAi_864,
       b4_nUAi_894,
       b4_nUAi_891,
       b4_nUAi_888,
       b4_nUAi_885,
       b4_nUAi_882,
       b4_nUAi_912,
       b4_nUAi_942,
       b4_nUAi_939,
       b4_nUAi_936,
       b4_nUAi_933,
       b4_nUAi_930,
       b4_nUAi_960,
       b4_nUAi_990,
       b4_nUAi_987,
       b4_nUAi_984,
       b4_nUAi_981,
       b4_nUAi_978,
       b4_nUAi_1008,
       b4_nUAi_1038,
       b4_nUAi_1035,
       b4_nUAi_1032,
       b4_nUAi_1029,
       b4_nUAi_1026,
       b4_nUAi_1056,
       b4_nUAi_1086,
       b4_nUAi_1083,
       b4_nUAi_1080,
       b4_nUAi_1077,
       b4_nUAi_1074,
       b4_nUAi_1107,
       b4_nUAi_1101,
       b4_nUAi_1095,
       b4_nUAi_1089,
       b6_2ZTGIf_6,
       b6_2ZTGIf_4,
       b6_2ZTGIf_3,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_7,
       b6_2ZTGIf_22,
       b6_2ZTGIf_20,
       b6_2ZTGIf_19,
       b6_2ZTGIf_18,
       b6_2ZTGIf_17,
       b6_2ZTGIf_16,
       b6_2ZTGIf_26,
       b6_2ZTGIf_25,
       b6_2ZTGIf_24,
       b6_2ZTGIf_23,
       b6_2ZTGIf_38,
       b6_2ZTGIf_36,
       b6_2ZTGIf_35,
       b6_2ZTGIf_34,
       b6_2ZTGIf_33,
       b6_2ZTGIf_32,
       b6_2ZTGIf_42,
       b6_2ZTGIf_41,
       b6_2ZTGIf_40,
       b6_2ZTGIf_39,
       b6_2ZTGIf_54,
       b6_2ZTGIf_52,
       b6_2ZTGIf_51,
       b6_2ZTGIf_50,
       b6_2ZTGIf_49,
       b6_2ZTGIf_48,
       b6_2ZTGIf_58,
       b6_2ZTGIf_57,
       b6_2ZTGIf_56,
       b6_2ZTGIf_55,
       b6_2ZTGIf_70,
       b6_2ZTGIf_68,
       b6_2ZTGIf_67,
       b6_2ZTGIf_66,
       b6_2ZTGIf_65,
       b6_2ZTGIf_64,
       b6_2ZTGIf_74,
       b6_2ZTGIf_73,
       b6_2ZTGIf_72,
       b6_2ZTGIf_71,
       b6_2ZTGIf_86,
       b6_2ZTGIf_84,
       b6_2ZTGIf_83,
       b6_2ZTGIf_82,
       b6_2ZTGIf_81,
       b6_2ZTGIf_80,
       b6_2ZTGIf_90,
       b6_2ZTGIf_89,
       b6_2ZTGIf_88,
       b6_2ZTGIf_87,
       b6_2ZTGIf_102,
       b6_2ZTGIf_100,
       b6_2ZTGIf_99,
       b6_2ZTGIf_98,
       b6_2ZTGIf_97,
       b6_2ZTGIf_96,
       b6_2ZTGIf_106,
       b6_2ZTGIf_105,
       b6_2ZTGIf_104,
       b6_2ZTGIf_103,
       b6_2ZTGIf_118,
       b6_2ZTGIf_116,
       b6_2ZTGIf_115,
       b6_2ZTGIf_114,
       b6_2ZTGIf_113,
       b6_2ZTGIf_112,
       b6_2ZTGIf_122,
       b6_2ZTGIf_121,
       b6_2ZTGIf_120,
       b6_2ZTGIf_119,
       b6_2ZTGIf_134,
       b6_2ZTGIf_132,
       b6_2ZTGIf_131,
       b6_2ZTGIf_130,
       b6_2ZTGIf_129,
       b6_2ZTGIf_128,
       b6_2ZTGIf_138,
       b6_2ZTGIf_137,
       b6_2ZTGIf_136,
       b6_2ZTGIf_135,
       b6_2ZTGIf_150,
       b6_2ZTGIf_148,
       b6_2ZTGIf_147,
       b6_2ZTGIf_146,
       b6_2ZTGIf_145,
       b6_2ZTGIf_144,
       b6_2ZTGIf_154,
       b6_2ZTGIf_153,
       b6_2ZTGIf_152,
       b6_2ZTGIf_151,
       b6_2ZTGIf_166,
       b6_2ZTGIf_164,
       b6_2ZTGIf_163,
       b6_2ZTGIf_162,
       b6_2ZTGIf_161,
       b6_2ZTGIf_160,
       b6_2ZTGIf_170,
       b6_2ZTGIf_169,
       b6_2ZTGIf_168,
       b6_2ZTGIf_167,
       b6_2ZTGIf_182,
       b6_2ZTGIf_180,
       b6_2ZTGIf_179,
       b6_2ZTGIf_178,
       b6_2ZTGIf_177,
       b6_2ZTGIf_176,
       b6_2ZTGIf_186,
       b6_2ZTGIf_185,
       b6_2ZTGIf_184,
       b6_2ZTGIf_183,
       b6_2ZTGIf_198,
       b6_2ZTGIf_196,
       b6_2ZTGIf_195,
       b6_2ZTGIf_194,
       b6_2ZTGIf_193,
       b6_2ZTGIf_192,
       b6_2ZTGIf_202,
       b6_2ZTGIf_201,
       b6_2ZTGIf_200,
       b6_2ZTGIf_199,
       b6_2ZTGIf_214,
       b6_2ZTGIf_212,
       b6_2ZTGIf_211,
       b6_2ZTGIf_210,
       b6_2ZTGIf_209,
       b6_2ZTGIf_208,
       b6_2ZTGIf_218,
       b6_2ZTGIf_217,
       b6_2ZTGIf_216,
       b6_2ZTGIf_215,
       b6_2ZTGIf_230,
       b6_2ZTGIf_228,
       b6_2ZTGIf_227,
       b6_2ZTGIf_226,
       b6_2ZTGIf_225,
       b6_2ZTGIf_224,
       b6_2ZTGIf_234,
       b6_2ZTGIf_233,
       b6_2ZTGIf_232,
       b6_2ZTGIf_231,
       b6_2ZTGIf_246,
       b6_2ZTGIf_244,
       b6_2ZTGIf_243,
       b6_2ZTGIf_242,
       b6_2ZTGIf_241,
       b6_2ZTGIf_240,
       b6_2ZTGIf_250,
       b6_2ZTGIf_249,
       b6_2ZTGIf_248,
       b6_2ZTGIf_247,
       b6_2ZTGIf_262,
       b6_2ZTGIf_260,
       b6_2ZTGIf_259,
       b6_2ZTGIf_258,
       b6_2ZTGIf_257,
       b6_2ZTGIf_256,
       b6_2ZTGIf_266,
       b6_2ZTGIf_265,
       b6_2ZTGIf_264,
       b6_2ZTGIf_263,
       b6_2ZTGIf_278,
       b6_2ZTGIf_276,
       b6_2ZTGIf_275,
       b6_2ZTGIf_274,
       b6_2ZTGIf_273,
       b6_2ZTGIf_272,
       b6_2ZTGIf_282,
       b6_2ZTGIf_281,
       b6_2ZTGIf_280,
       b6_2ZTGIf_279,
       b6_2ZTGIf_294,
       b6_2ZTGIf_292,
       b6_2ZTGIf_291,
       b6_2ZTGIf_290,
       b6_2ZTGIf_289,
       b6_2ZTGIf_288,
       b6_2ZTGIf_298,
       b6_2ZTGIf_297,
       b6_2ZTGIf_296,
       b6_2ZTGIf_295,
       b6_2ZTGIf_310,
       b6_2ZTGIf_308,
       b6_2ZTGIf_307,
       b6_2ZTGIf_306,
       b6_2ZTGIf_305,
       b6_2ZTGIf_304,
       b6_2ZTGIf_314,
       b6_2ZTGIf_313,
       b6_2ZTGIf_312,
       b6_2ZTGIf_311,
       b6_2ZTGIf_326,
       b6_2ZTGIf_324,
       b6_2ZTGIf_323,
       b6_2ZTGIf_322,
       b6_2ZTGIf_321,
       b6_2ZTGIf_320,
       b6_2ZTGIf_330,
       b6_2ZTGIf_329,
       b6_2ZTGIf_328,
       b6_2ZTGIf_327,
       b6_2ZTGIf_342,
       b6_2ZTGIf_340,
       b6_2ZTGIf_339,
       b6_2ZTGIf_338,
       b6_2ZTGIf_337,
       b6_2ZTGIf_336,
       b6_2ZTGIf_346,
       b6_2ZTGIf_345,
       b6_2ZTGIf_344,
       b6_2ZTGIf_343,
       b6_2ZTGIf_358,
       b6_2ZTGIf_356,
       b6_2ZTGIf_355,
       b6_2ZTGIf_354,
       b6_2ZTGIf_353,
       b6_2ZTGIf_352,
       b6_2ZTGIf_362,
       b6_2ZTGIf_361,
       b6_2ZTGIf_360,
       b6_2ZTGIf_359,
       b6_2ZTGIf_375,
       b6_2ZTGIf_373,
       b6_2ZTGIf_371,
       b6_2ZTGIf_369,
       BW_clk_c,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4,
       N_25_5,
       N_27_5,
       N_25_6,
       N_27_6,
       N_25_7,
       N_27_7,
       N_25_8,
       N_27_8,
       N_25_9,
       N_27_9,
       N_25_10,
       N_27_10,
       N_25_11,
       N_27_11,
       N_25_12,
       N_27_12,
       N_25_13,
       N_27_13,
       N_25_14,
       N_27_14,
       N_25_15,
       N_27_15,
       N_25_16,
       N_27_16,
       N_25_17,
       N_27_17,
       N_25_18,
       N_27_18,
       N_25_19,
       N_27_19,
       N_25_20,
       N_27_20,
       N_25_21,
       N_27_21,
       N_25_22,
       N_27_22,
       N_25_23,
       N_27_23,
       N_25_24,
       N_27_24,
       N_25_25,
       N_27_25,
       N_25_26,
       N_27_26,
       N_25_27,
       N_27_27,
       N_25_28,
       N_27_28,
       N_25_29,
       N_27_29,
       N_25_30,
       N_27_30,
       N_25_31,
       N_27_31,
       N_25_32,
       N_27_32,
       N_25_33,
       N_27_33,
       N_25_34,
       N_27_34,
       N_25_35,
       N_27_35,
       N_25_36,
       N_27_36,
       N_25_37,
       N_27_37,
       N_25_38,
       N_27_38,
       N_25_39,
       N_27_39,
       N_25_40,
       N_27_40,
       N_25_41,
       N_27_41,
       N_25_42,
       N_27_42,
       N_25_43,
       N_27_43,
       N_25_44,
       N_27_44,
       N_25_45,
       N_27_45,
       N_25_46,
       N_27_46,
       N_25_47,
       N_27_47,
       N_25_48,
       N_27_48,
       N_25_49,
       N_27_49,
       N_25_50,
       N_27_50,
       N_25_51,
       N_27_51,
       N_25_52,
       N_27_52,
       N_25_53,
       N_27_53,
       N_25_54,
       N_27_54,
       N_25_55,
       N_27_55,
       N_25_56,
       N_27_56,
       N_25_57,
       N_27_57,
       N_25_58,
       N_27_58,
       N_25_59,
       N_27_59,
       N_25_60,
       N_27_60,
       N_25_61,
       N_27_61,
       N_25_62,
       N_27_62,
       N_25_63,
       N_27_63,
       N_25_64,
       N_27_64,
       N_25_65,
       N_27_65,
       N_25_66,
       N_27_66,
       N_25_67,
       N_27_67,
       N_25_68,
       N_27_68,
       N_25_69,
       N_27_69,
       N_25_70,
       N_27_70,
       N_25_71,
       N_27_71,
       N_25_72,
       N_27_72,
       N_25_73,
       N_27_73,
       N_25_74,
       N_27_74,
       N_25_75,
       N_27_75,
       N_25_76,
       N_27_76,
       N_25_77,
       N_27_77,
       N_25_78,
       N_27_78,
       N_25_79,
       N_27_79,
       N_25_80,
       N_27_80,
       N_25_81,
       N_27_81,
       N_25_82,
       N_27_82,
       N_25_83,
       N_27_83,
       N_25_84,
       N_27_84,
       N_25_85,
       N_27_85,
       N_25_86,
       N_27_86,
       N_25_87,
       N_27_87,
       N_25_88,
       N_27_88,
       N_25_89,
       N_27_89,
       N_25_90,
       N_27_90,
       N_25_91,
       N_27_91,
       N_25_92,
       N_27_92,
       N_25_93,
       N_27_93,
       N_25_94,
       N_27_94,
       N_25_95,
       N_27_95,
       N_25_96,
       N_27_96,
       N_25_97,
       N_27_97,
       N_25_98,
       N_27_98,
       N_25_99,
       N_27_99,
       N_25_100,
       N_27_100,
       N_25_101,
       N_27_101,
       N_25_102,
       N_27_102,
       N_25_103,
       N_27_103,
       N_25_104,
       N_27_104,
       N_25_105,
       N_27_105,
       N_25_106,
       N_27_106,
       N_25_107,
       N_27_107,
       N_25_108,
       N_27_108,
       N_25_109,
       N_27_109,
       N_25_110,
       N_27_110,
       N_25_111,
       N_27_111,
       N_25_112,
       N_27_112,
       N_25_113,
       N_27_113,
       N_25_114,
       N_27_114,
       N_25_115,
       N_27_115,
       N_25_116,
       N_27_116,
       N_25_117,
       N_27_117,
       N_25_118,
       N_27_118,
       N_25_119,
       N_27_119,
       N_25_120,
       N_27_120,
       N_25_121,
       N_27_121,
       N_25_122,
       N_27_122,
       N_25_123,
       N_27_123,
       N_25_124,
       N_27_124,
       N_25_125,
       N_27_125,
       N_25_126,
       N_27_126,
       N_25_127,
       N_27_127,
       N_25_128,
       N_27_128,
       N_25_129,
       N_27_129,
       N_25_130,
       N_27_130,
       N_25_131,
       N_27_131,
       N_25_132,
       N_27_132,
       N_25_133,
       N_27_133,
       N_25_134,
       N_27_134,
       N_25_135,
       N_27_135,
       N_25_136,
       N_27_136,
       N_25_137,
       N_27_137,
       N_25_138,
       N_27_138,
       N_25_139,
       N_27_139,
       N_25_140,
       N_27_140,
       N_25_141,
       b7_PSyi3wy,
       N_27_141
    );
output [1:1] b11_uUT0JC4gFrY;
input  b4_nUAi_0;
input  b4_nUAi_30;
input  b4_nUAi_27;
input  b4_nUAi_24;
input  b4_nUAi_21;
input  b4_nUAi_18;
input  b4_nUAi_48;
input  b4_nUAi_78;
input  b4_nUAi_75;
input  b4_nUAi_72;
input  b4_nUAi_69;
input  b4_nUAi_66;
input  b4_nUAi_96;
input  b4_nUAi_126;
input  b4_nUAi_123;
input  b4_nUAi_120;
input  b4_nUAi_117;
input  b4_nUAi_114;
input  b4_nUAi_144;
input  b4_nUAi_174;
input  b4_nUAi_171;
input  b4_nUAi_168;
input  b4_nUAi_165;
input  b4_nUAi_162;
input  b4_nUAi_192;
input  b4_nUAi_222;
input  b4_nUAi_219;
input  b4_nUAi_216;
input  b4_nUAi_213;
input  b4_nUAi_210;
input  b4_nUAi_240;
input  b4_nUAi_270;
input  b4_nUAi_267;
input  b4_nUAi_264;
input  b4_nUAi_261;
input  b4_nUAi_258;
input  b4_nUAi_288;
input  b4_nUAi_318;
input  b4_nUAi_315;
input  b4_nUAi_312;
input  b4_nUAi_309;
input  b4_nUAi_306;
input  b4_nUAi_336;
input  b4_nUAi_366;
input  b4_nUAi_363;
input  b4_nUAi_360;
input  b4_nUAi_357;
input  b4_nUAi_354;
input  b4_nUAi_384;
input  b4_nUAi_414;
input  b4_nUAi_411;
input  b4_nUAi_408;
input  b4_nUAi_405;
input  b4_nUAi_402;
input  b4_nUAi_432;
input  b4_nUAi_462;
input  b4_nUAi_459;
input  b4_nUAi_456;
input  b4_nUAi_453;
input  b4_nUAi_450;
input  b4_nUAi_480;
input  b4_nUAi_510;
input  b4_nUAi_507;
input  b4_nUAi_504;
input  b4_nUAi_501;
input  b4_nUAi_498;
input  b4_nUAi_528;
input  b4_nUAi_558;
input  b4_nUAi_555;
input  b4_nUAi_552;
input  b4_nUAi_549;
input  b4_nUAi_546;
input  b4_nUAi_576;
input  b4_nUAi_606;
input  b4_nUAi_603;
input  b4_nUAi_600;
input  b4_nUAi_597;
input  b4_nUAi_594;
input  b4_nUAi_624;
input  b4_nUAi_654;
input  b4_nUAi_651;
input  b4_nUAi_648;
input  b4_nUAi_645;
input  b4_nUAi_642;
input  b4_nUAi_672;
input  b4_nUAi_702;
input  b4_nUAi_699;
input  b4_nUAi_696;
input  b4_nUAi_693;
input  b4_nUAi_690;
input  b4_nUAi_720;
input  b4_nUAi_750;
input  b4_nUAi_747;
input  b4_nUAi_744;
input  b4_nUAi_741;
input  b4_nUAi_738;
input  b4_nUAi_768;
input  b4_nUAi_798;
input  b4_nUAi_795;
input  b4_nUAi_792;
input  b4_nUAi_789;
input  b4_nUAi_786;
input  b4_nUAi_816;
input  b4_nUAi_846;
input  b4_nUAi_843;
input  b4_nUAi_840;
input  b4_nUAi_837;
input  b4_nUAi_834;
input  b4_nUAi_864;
input  b4_nUAi_894;
input  b4_nUAi_891;
input  b4_nUAi_888;
input  b4_nUAi_885;
input  b4_nUAi_882;
input  b4_nUAi_912;
input  b4_nUAi_942;
input  b4_nUAi_939;
input  b4_nUAi_936;
input  b4_nUAi_933;
input  b4_nUAi_930;
input  b4_nUAi_960;
input  b4_nUAi_990;
input  b4_nUAi_987;
input  b4_nUAi_984;
input  b4_nUAi_981;
input  b4_nUAi_978;
input  b4_nUAi_1008;
input  b4_nUAi_1038;
input  b4_nUAi_1035;
input  b4_nUAi_1032;
input  b4_nUAi_1029;
input  b4_nUAi_1026;
input  b4_nUAi_1056;
input  b4_nUAi_1086;
input  b4_nUAi_1083;
input  b4_nUAi_1080;
input  b4_nUAi_1077;
input  b4_nUAi_1074;
input  b4_nUAi_1107;
input  b4_nUAi_1101;
input  b4_nUAi_1095;
input  b4_nUAi_1089;
input  b6_2ZTGIf_6;
input  b6_2ZTGIf_4;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_22;
input  b6_2ZTGIf_20;
input  b6_2ZTGIf_19;
input  b6_2ZTGIf_18;
input  b6_2ZTGIf_17;
input  b6_2ZTGIf_16;
input  b6_2ZTGIf_26;
input  b6_2ZTGIf_25;
input  b6_2ZTGIf_24;
input  b6_2ZTGIf_23;
input  b6_2ZTGIf_38;
input  b6_2ZTGIf_36;
input  b6_2ZTGIf_35;
input  b6_2ZTGIf_34;
input  b6_2ZTGIf_33;
input  b6_2ZTGIf_32;
input  b6_2ZTGIf_42;
input  b6_2ZTGIf_41;
input  b6_2ZTGIf_40;
input  b6_2ZTGIf_39;
input  b6_2ZTGIf_54;
input  b6_2ZTGIf_52;
input  b6_2ZTGIf_51;
input  b6_2ZTGIf_50;
input  b6_2ZTGIf_49;
input  b6_2ZTGIf_48;
input  b6_2ZTGIf_58;
input  b6_2ZTGIf_57;
input  b6_2ZTGIf_56;
input  b6_2ZTGIf_55;
input  b6_2ZTGIf_70;
input  b6_2ZTGIf_68;
input  b6_2ZTGIf_67;
input  b6_2ZTGIf_66;
input  b6_2ZTGIf_65;
input  b6_2ZTGIf_64;
input  b6_2ZTGIf_74;
input  b6_2ZTGIf_73;
input  b6_2ZTGIf_72;
input  b6_2ZTGIf_71;
input  b6_2ZTGIf_86;
input  b6_2ZTGIf_84;
input  b6_2ZTGIf_83;
input  b6_2ZTGIf_82;
input  b6_2ZTGIf_81;
input  b6_2ZTGIf_80;
input  b6_2ZTGIf_90;
input  b6_2ZTGIf_89;
input  b6_2ZTGIf_88;
input  b6_2ZTGIf_87;
input  b6_2ZTGIf_102;
input  b6_2ZTGIf_100;
input  b6_2ZTGIf_99;
input  b6_2ZTGIf_98;
input  b6_2ZTGIf_97;
input  b6_2ZTGIf_96;
input  b6_2ZTGIf_106;
input  b6_2ZTGIf_105;
input  b6_2ZTGIf_104;
input  b6_2ZTGIf_103;
input  b6_2ZTGIf_118;
input  b6_2ZTGIf_116;
input  b6_2ZTGIf_115;
input  b6_2ZTGIf_114;
input  b6_2ZTGIf_113;
input  b6_2ZTGIf_112;
input  b6_2ZTGIf_122;
input  b6_2ZTGIf_121;
input  b6_2ZTGIf_120;
input  b6_2ZTGIf_119;
input  b6_2ZTGIf_134;
input  b6_2ZTGIf_132;
input  b6_2ZTGIf_131;
input  b6_2ZTGIf_130;
input  b6_2ZTGIf_129;
input  b6_2ZTGIf_128;
input  b6_2ZTGIf_138;
input  b6_2ZTGIf_137;
input  b6_2ZTGIf_136;
input  b6_2ZTGIf_135;
input  b6_2ZTGIf_150;
input  b6_2ZTGIf_148;
input  b6_2ZTGIf_147;
input  b6_2ZTGIf_146;
input  b6_2ZTGIf_145;
input  b6_2ZTGIf_144;
input  b6_2ZTGIf_154;
input  b6_2ZTGIf_153;
input  b6_2ZTGIf_152;
input  b6_2ZTGIf_151;
input  b6_2ZTGIf_166;
input  b6_2ZTGIf_164;
input  b6_2ZTGIf_163;
input  b6_2ZTGIf_162;
input  b6_2ZTGIf_161;
input  b6_2ZTGIf_160;
input  b6_2ZTGIf_170;
input  b6_2ZTGIf_169;
input  b6_2ZTGIf_168;
input  b6_2ZTGIf_167;
input  b6_2ZTGIf_182;
input  b6_2ZTGIf_180;
input  b6_2ZTGIf_179;
input  b6_2ZTGIf_178;
input  b6_2ZTGIf_177;
input  b6_2ZTGIf_176;
input  b6_2ZTGIf_186;
input  b6_2ZTGIf_185;
input  b6_2ZTGIf_184;
input  b6_2ZTGIf_183;
input  b6_2ZTGIf_198;
input  b6_2ZTGIf_196;
input  b6_2ZTGIf_195;
input  b6_2ZTGIf_194;
input  b6_2ZTGIf_193;
input  b6_2ZTGIf_192;
input  b6_2ZTGIf_202;
input  b6_2ZTGIf_201;
input  b6_2ZTGIf_200;
input  b6_2ZTGIf_199;
input  b6_2ZTGIf_214;
input  b6_2ZTGIf_212;
input  b6_2ZTGIf_211;
input  b6_2ZTGIf_210;
input  b6_2ZTGIf_209;
input  b6_2ZTGIf_208;
input  b6_2ZTGIf_218;
input  b6_2ZTGIf_217;
input  b6_2ZTGIf_216;
input  b6_2ZTGIf_215;
input  b6_2ZTGIf_230;
input  b6_2ZTGIf_228;
input  b6_2ZTGIf_227;
input  b6_2ZTGIf_226;
input  b6_2ZTGIf_225;
input  b6_2ZTGIf_224;
input  b6_2ZTGIf_234;
input  b6_2ZTGIf_233;
input  b6_2ZTGIf_232;
input  b6_2ZTGIf_231;
input  b6_2ZTGIf_246;
input  b6_2ZTGIf_244;
input  b6_2ZTGIf_243;
input  b6_2ZTGIf_242;
input  b6_2ZTGIf_241;
input  b6_2ZTGIf_240;
input  b6_2ZTGIf_250;
input  b6_2ZTGIf_249;
input  b6_2ZTGIf_248;
input  b6_2ZTGIf_247;
input  b6_2ZTGIf_262;
input  b6_2ZTGIf_260;
input  b6_2ZTGIf_259;
input  b6_2ZTGIf_258;
input  b6_2ZTGIf_257;
input  b6_2ZTGIf_256;
input  b6_2ZTGIf_266;
input  b6_2ZTGIf_265;
input  b6_2ZTGIf_264;
input  b6_2ZTGIf_263;
input  b6_2ZTGIf_278;
input  b6_2ZTGIf_276;
input  b6_2ZTGIf_275;
input  b6_2ZTGIf_274;
input  b6_2ZTGIf_273;
input  b6_2ZTGIf_272;
input  b6_2ZTGIf_282;
input  b6_2ZTGIf_281;
input  b6_2ZTGIf_280;
input  b6_2ZTGIf_279;
input  b6_2ZTGIf_294;
input  b6_2ZTGIf_292;
input  b6_2ZTGIf_291;
input  b6_2ZTGIf_290;
input  b6_2ZTGIf_289;
input  b6_2ZTGIf_288;
input  b6_2ZTGIf_298;
input  b6_2ZTGIf_297;
input  b6_2ZTGIf_296;
input  b6_2ZTGIf_295;
input  b6_2ZTGIf_310;
input  b6_2ZTGIf_308;
input  b6_2ZTGIf_307;
input  b6_2ZTGIf_306;
input  b6_2ZTGIf_305;
input  b6_2ZTGIf_304;
input  b6_2ZTGIf_314;
input  b6_2ZTGIf_313;
input  b6_2ZTGIf_312;
input  b6_2ZTGIf_311;
input  b6_2ZTGIf_326;
input  b6_2ZTGIf_324;
input  b6_2ZTGIf_323;
input  b6_2ZTGIf_322;
input  b6_2ZTGIf_321;
input  b6_2ZTGIf_320;
input  b6_2ZTGIf_330;
input  b6_2ZTGIf_329;
input  b6_2ZTGIf_328;
input  b6_2ZTGIf_327;
input  b6_2ZTGIf_342;
input  b6_2ZTGIf_340;
input  b6_2ZTGIf_339;
input  b6_2ZTGIf_338;
input  b6_2ZTGIf_337;
input  b6_2ZTGIf_336;
input  b6_2ZTGIf_346;
input  b6_2ZTGIf_345;
input  b6_2ZTGIf_344;
input  b6_2ZTGIf_343;
input  b6_2ZTGIf_358;
input  b6_2ZTGIf_356;
input  b6_2ZTGIf_355;
input  b6_2ZTGIf_354;
input  b6_2ZTGIf_353;
input  b6_2ZTGIf_352;
input  b6_2ZTGIf_362;
input  b6_2ZTGIf_361;
input  b6_2ZTGIf_360;
input  b6_2ZTGIf_359;
input  b6_2ZTGIf_375;
input  b6_2ZTGIf_373;
input  b6_2ZTGIf_371;
input  b6_2ZTGIf_369;
input  BW_clk_c;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;
input  N_25_5;
input  N_27_5;
input  N_25_6;
input  N_27_6;
input  N_25_7;
input  N_27_7;
input  N_25_8;
input  N_27_8;
input  N_25_9;
input  N_27_9;
input  N_25_10;
input  N_27_10;
input  N_25_11;
input  N_27_11;
input  N_25_12;
input  N_27_12;
input  N_25_13;
input  N_27_13;
input  N_25_14;
input  N_27_14;
input  N_25_15;
input  N_27_15;
input  N_25_16;
input  N_27_16;
input  N_25_17;
input  N_27_17;
input  N_25_18;
input  N_27_18;
input  N_25_19;
input  N_27_19;
input  N_25_20;
input  N_27_20;
input  N_25_21;
input  N_27_21;
input  N_25_22;
input  N_27_22;
input  N_25_23;
input  N_27_23;
input  N_25_24;
input  N_27_24;
input  N_25_25;
input  N_27_25;
input  N_25_26;
input  N_27_26;
input  N_25_27;
input  N_27_27;
input  N_25_28;
input  N_27_28;
input  N_25_29;
input  N_27_29;
input  N_25_30;
input  N_27_30;
input  N_25_31;
input  N_27_31;
input  N_25_32;
input  N_27_32;
input  N_25_33;
input  N_27_33;
input  N_25_34;
input  N_27_34;
input  N_25_35;
input  N_27_35;
input  N_25_36;
input  N_27_36;
input  N_25_37;
input  N_27_37;
input  N_25_38;
input  N_27_38;
input  N_25_39;
input  N_27_39;
input  N_25_40;
input  N_27_40;
input  N_25_41;
input  N_27_41;
input  N_25_42;
input  N_27_42;
input  N_25_43;
input  N_27_43;
input  N_25_44;
input  N_27_44;
input  N_25_45;
input  N_27_45;
input  N_25_46;
input  N_27_46;
input  N_25_47;
input  N_27_47;
input  N_25_48;
input  N_27_48;
input  N_25_49;
input  N_27_49;
input  N_25_50;
input  N_27_50;
input  N_25_51;
input  N_27_51;
input  N_25_52;
input  N_27_52;
input  N_25_53;
input  N_27_53;
input  N_25_54;
input  N_27_54;
input  N_25_55;
input  N_27_55;
input  N_25_56;
input  N_27_56;
input  N_25_57;
input  N_27_57;
input  N_25_58;
input  N_27_58;
input  N_25_59;
input  N_27_59;
input  N_25_60;
input  N_27_60;
input  N_25_61;
input  N_27_61;
input  N_25_62;
input  N_27_62;
input  N_25_63;
input  N_27_63;
input  N_25_64;
input  N_27_64;
input  N_25_65;
input  N_27_65;
input  N_25_66;
input  N_27_66;
input  N_25_67;
input  N_27_67;
input  N_25_68;
input  N_27_68;
input  N_25_69;
input  N_27_69;
input  N_25_70;
input  N_27_70;
input  N_25_71;
input  N_27_71;
input  N_25_72;
input  N_27_72;
input  N_25_73;
input  N_27_73;
input  N_25_74;
input  N_27_74;
input  N_25_75;
input  N_27_75;
input  N_25_76;
input  N_27_76;
input  N_25_77;
input  N_27_77;
input  N_25_78;
input  N_27_78;
input  N_25_79;
input  N_27_79;
input  N_25_80;
input  N_27_80;
input  N_25_81;
input  N_27_81;
input  N_25_82;
input  N_27_82;
input  N_25_83;
input  N_27_83;
input  N_25_84;
input  N_27_84;
input  N_25_85;
input  N_27_85;
input  N_25_86;
input  N_27_86;
input  N_25_87;
input  N_27_87;
input  N_25_88;
input  N_27_88;
input  N_25_89;
input  N_27_89;
input  N_25_90;
input  N_27_90;
input  N_25_91;
input  N_27_91;
input  N_25_92;
input  N_27_92;
input  N_25_93;
input  N_27_93;
input  N_25_94;
input  N_27_94;
input  N_25_95;
input  N_27_95;
input  N_25_96;
input  N_27_96;
input  N_25_97;
input  N_27_97;
input  N_25_98;
input  N_27_98;
input  N_25_99;
input  N_27_99;
input  N_25_100;
input  N_27_100;
input  N_25_101;
input  N_27_101;
input  N_25_102;
input  N_27_102;
input  N_25_103;
input  N_27_103;
input  N_25_104;
input  N_27_104;
input  N_25_105;
input  N_27_105;
input  N_25_106;
input  N_27_106;
input  N_25_107;
input  N_27_107;
input  N_25_108;
input  N_27_108;
input  N_25_109;
input  N_27_109;
input  N_25_110;
input  N_27_110;
input  N_25_111;
input  N_27_111;
input  N_25_112;
input  N_27_112;
input  N_25_113;
input  N_27_113;
input  N_25_114;
input  N_27_114;
input  N_25_115;
input  N_27_115;
input  N_25_116;
input  N_27_116;
input  N_25_117;
input  N_27_117;
input  N_25_118;
input  N_27_118;
input  N_25_119;
input  N_27_119;
input  N_25_120;
input  N_27_120;
input  N_25_121;
input  N_27_121;
input  N_25_122;
input  N_27_122;
input  N_25_123;
input  N_27_123;
input  N_25_124;
input  N_27_124;
input  N_25_125;
input  N_27_125;
input  N_25_126;
input  N_27_126;
input  N_25_127;
input  N_27_127;
input  N_25_128;
input  N_27_128;
input  N_25_129;
input  N_27_129;
input  N_25_130;
input  N_27_130;
input  N_25_131;
input  N_27_131;
input  N_25_132;
input  N_27_132;
input  N_25_133;
input  N_27_133;
input  N_25_134;
input  N_27_134;
input  N_25_135;
input  N_27_135;
input  N_25_136;
input  N_27_136;
input  N_25_137;
input  N_27_137;
input  N_25_138;
input  N_27_138;
input  N_25_139;
input  N_27_139;
input  N_25_140;
input  N_27_140;
input  N_25_141;
input  b7_PSyi3wy;
input  N_27_141;

    wire \b14_CZS0wfY_d_FH9m[7]_net_1 , VCC_net_1, 
        \b13_CZS0wfY_d_FH9[7] , GND_net_1, 
        \b14_CZS0wfY_d_FH9m[6]_net_1 , \b13_CZS0wfY_d_FH9[6] , 
        \b14_CZS0wfY_d_FH9m[5]_net_1 , \b13_CZS0wfY_d_FH9[5] , 
        \b14_CZS0wfY_d_FH9m[4]_net_1 , \b13_CZS0wfY_d_FH9[4] , 
        \b14_CZS0wfY_d_FH9m[3]_net_1 , \b13_CZS0wfY_d_FH9[3] , 
        \b14_CZS0wfY_d_FH9m[2]_net_1 , \b13_CZS0wfY_d_FH9[2] , 
        \b14_CZS0wfY_d_FH9m[1]_net_1 , \b13_CZS0wfY_d_FH9[1] , 
        \b14_CZS0wfY_d_FH9m[0]_net_1 , \b13_CZS0wfY_d_FH9[0] , 
        \b14_CZS0wfY_d_FH9m[22]_net_1 , \b13_CZS0wfY_d_FH9[22] , 
        \b14_CZS0wfY_d_FH9m[21]_net_1 , \b13_CZS0wfY_d_FH9[21] , 
        \b14_CZS0wfY_d_FH9m[20]_net_1 , \b13_CZS0wfY_d_FH9[20] , 
        \b14_CZS0wfY_d_FH9m[19]_net_1 , \b13_CZS0wfY_d_FH9[19] , 
        \b14_CZS0wfY_d_FH9m[18]_net_1 , \b13_CZS0wfY_d_FH9[18] , 
        \b14_CZS0wfY_d_FH9m[17]_net_1 , \b13_CZS0wfY_d_FH9[17] , 
        \b14_CZS0wfY_d_FH9m[16]_net_1 , \b13_CZS0wfY_d_FH9[16] , 
        \b14_CZS0wfY_d_FH9m[15]_net_1 , \b13_CZS0wfY_d_FH9[15] , 
        \b14_CZS0wfY_d_FH9m[14]_net_1 , \b13_CZS0wfY_d_FH9[14] , 
        \b14_CZS0wfY_d_FH9m[13]_net_1 , \b13_CZS0wfY_d_FH9[13] , 
        \b14_CZS0wfY_d_FH9m[12]_net_1 , \b13_CZS0wfY_d_FH9[12] , 
        \b14_CZS0wfY_d_FH9m[11]_net_1 , \b13_CZS0wfY_d_FH9[11] , 
        \b14_CZS0wfY_d_FH9m[10]_net_1 , \b13_CZS0wfY_d_FH9[10] , 
        \b14_CZS0wfY_d_FH9m[9]_net_1 , \b13_CZS0wfY_d_FH9[9] , 
        \b14_CZS0wfY_d_FH9m[8]_net_1 , \b13_CZS0wfY_d_FH9[8] , 
        \b14_CZS0wfY_d_FH9m[23]_net_1 , \b13_CZS0wfY_d_FH9[23] ;
    
    b9_O2yyf_fG2_x_22_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_a6 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[10] }), .b4_nUAi_0(
        b4_nUAi_480), .b4_nUAi_30(b4_nUAi_510), .b4_nUAi_27(
        b4_nUAi_507), .b4_nUAi_24(b4_nUAi_504), .b4_nUAi_21(
        b4_nUAi_501), .b4_nUAi_18(b4_nUAi_498), .b6_2ZTGIf_6(
        b6_2ZTGIf_166), .b6_2ZTGIf_4(b6_2ZTGIf_164), .b6_2ZTGIf_3(
        b6_2ZTGIf_163), .b6_2ZTGIf_2(b6_2ZTGIf_162), .b6_2ZTGIf_1(
        b6_2ZTGIf_161), .b6_2ZTGIf_0(b6_2ZTGIf_160), .b6_2ZTGIf_10(
        b6_2ZTGIf_170), .b6_2ZTGIf_9(b6_2ZTGIf_169), .b6_2ZTGIf_8(
        b6_2ZTGIf_168), .b6_2ZTGIf_7(b6_2ZTGIf_167), .N_25(N_25_59), 
        .N_27(N_27_59), .N_25_0(N_25_60), .N_27_0(N_27_60), .N_25_1(
        N_25_61), .N_27_1(N_27_61), .N_25_2(N_25_62), .N_27_2(N_27_62), 
        .N_25_3(N_25_63), .N_27_3(N_27_63), .N_25_4(N_25_64), .N_27_4(
        N_27_64));
    b9_O2yyf_fG2_x_17_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_a9 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[15] }), .b4_nUAi_0(
        b4_nUAi_720), .b4_nUAi_30(b4_nUAi_750), .b4_nUAi_27(
        b4_nUAi_747), .b4_nUAi_24(b4_nUAi_744), .b4_nUAi_21(
        b4_nUAi_741), .b4_nUAi_18(b4_nUAi_738), .b6_2ZTGIf_6(
        b6_2ZTGIf_246), .b6_2ZTGIf_4(b6_2ZTGIf_244), .b6_2ZTGIf_3(
        b6_2ZTGIf_243), .b6_2ZTGIf_2(b6_2ZTGIf_242), .b6_2ZTGIf_1(
        b6_2ZTGIf_241), .b6_2ZTGIf_0(b6_2ZTGIf_240), .b6_2ZTGIf_10(
        b6_2ZTGIf_250), .b6_2ZTGIf_9(b6_2ZTGIf_249), .b6_2ZTGIf_8(
        b6_2ZTGIf_248), .b6_2ZTGIf_7(b6_2ZTGIf_247), .N_25(N_25_89), 
        .N_27(N_27_89), .N_25_0(N_25_90), .N_27_0(N_27_90), .N_25_1(
        N_25_91), .N_27_1(N_27_91), .N_25_2(N_25_92), .N_27_2(N_27_92), 
        .N_25_3(N_25_93), .N_27_3(N_27_93), .N_25_4(N_25_94), .N_27_4(
        N_27_94));
    b9_O2yyf_fG2_x_14_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_aC (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[18] }), .b4_nUAi_0(
        b4_nUAi_864), .b4_nUAi_30(b4_nUAi_894), .b4_nUAi_27(
        b4_nUAi_891), .b4_nUAi_24(b4_nUAi_888), .b4_nUAi_21(
        b4_nUAi_885), .b4_nUAi_18(b4_nUAi_882), .b6_2ZTGIf_6(
        b6_2ZTGIf_294), .b6_2ZTGIf_4(b6_2ZTGIf_292), .b6_2ZTGIf_3(
        b6_2ZTGIf_291), .b6_2ZTGIf_2(b6_2ZTGIf_290), .b6_2ZTGIf_1(
        b6_2ZTGIf_289), .b6_2ZTGIf_0(b6_2ZTGIf_288), .b6_2ZTGIf_10(
        b6_2ZTGIf_298), .b6_2ZTGIf_9(b6_2ZTGIf_297), .b6_2ZTGIf_8(
        b6_2ZTGIf_296), .b6_2ZTGIf_7(b6_2ZTGIf_295), .N_25(N_25_107), 
        .N_27(N_27_107), .N_25_0(N_25_108), .N_27_0(N_27_108), .N_25_1(
        N_25_109), .N_27_1(N_27_109), .N_25_2(N_25_110), .N_27_2(
        N_27_110), .N_25_3(N_25_111), .N_27_3(N_27_111), .N_25_4(
        N_25_112), .N_27_4(N_27_112));
    b9_O2yyf_fG2_x_29_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_I (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[3] }), .b4_nUAi_0(
        b4_nUAi_144), .b4_nUAi_30(b4_nUAi_174), .b4_nUAi_27(
        b4_nUAi_171), .b4_nUAi_24(b4_nUAi_168), .b4_nUAi_21(
        b4_nUAi_165), .b4_nUAi_18(b4_nUAi_162), .b6_2ZTGIf_6(
        b6_2ZTGIf_54), .b6_2ZTGIf_4(b6_2ZTGIf_52), .b6_2ZTGIf_3(
        b6_2ZTGIf_51), .b6_2ZTGIf_2(b6_2ZTGIf_50), .b6_2ZTGIf_1(
        b6_2ZTGIf_49), .b6_2ZTGIf_0(b6_2ZTGIf_48), .b6_2ZTGIf_10(
        b6_2ZTGIf_58), .b6_2ZTGIf_9(b6_2ZTGIf_57), .b6_2ZTGIf_8(
        b6_2ZTGIf_56), .b6_2ZTGIf_7(b6_2ZTGIf_55), .N_25(N_25_17), 
        .N_27(N_27_17), .N_25_0(N_25_18), .N_27_0(N_27_18), .N_25_1(
        N_25_19), .N_27_1(N_27_19), .N_25_2(N_25_20), .N_27_2(N_27_20), 
        .N_25_3(N_25_21), .N_27_3(N_27_21), .N_25_4(N_25_22), .N_27_4(
        N_27_22));
    SLE \b14_CZS0wfY_d_FH9m[15]  (.D(\b13_CZS0wfY_d_FH9[15] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[15]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[3]  (.D(\b13_CZS0wfY_d_FH9[3] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[3]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[10]  (.D(\b13_CZS0wfY_d_FH9[10] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[10]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[19]  (.D(\b13_CZS0wfY_d_FH9[19] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[19]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[17]  (.D(\b13_CZS0wfY_d_FH9[17] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[17]_net_1 ));
    b9_O2yyf_fG2_x_19_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_aF (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[13] }), .b4_nUAi_0(
        b4_nUAi_624), .b4_nUAi_30(b4_nUAi_654), .b4_nUAi_27(
        b4_nUAi_651), .b4_nUAi_24(b4_nUAi_648), .b4_nUAi_21(
        b4_nUAi_645), .b4_nUAi_18(b4_nUAi_642), .b6_2ZTGIf_6(
        b6_2ZTGIf_214), .b6_2ZTGIf_4(b6_2ZTGIf_212), .b6_2ZTGIf_3(
        b6_2ZTGIf_211), .b6_2ZTGIf_2(b6_2ZTGIf_210), .b6_2ZTGIf_1(
        b6_2ZTGIf_209), .b6_2ZTGIf_0(b6_2ZTGIf_208), .b6_2ZTGIf_10(
        b6_2ZTGIf_218), .b6_2ZTGIf_9(b6_2ZTGIf_217), .b6_2ZTGIf_8(
        b6_2ZTGIf_216), .b6_2ZTGIf_7(b6_2ZTGIf_215), .N_25(N_25_77), 
        .N_27(N_27_77), .N_25_0(N_25_78), .N_27_0(N_27_78), .N_25_1(
        N_25_79), .N_27_1(N_27_79), .N_25_2(N_25_80), .N_27_2(N_27_80), 
        .N_25_3(N_25_81), .N_27_3(N_27_81), .N_25_4(N_25_82), .N_27_4(
        N_27_82));
    SLE \b14_CZS0wfY_d_FH9m[7]  (.D(\b13_CZS0wfY_d_FH9[7] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[7]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[12]  (.D(\b13_CZS0wfY_d_FH9[12] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[12]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[23]  (.D(\b13_CZS0wfY_d_FH9[23] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[23]_net_1 ));
    b9_O2yyf_fG2_x_26_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_S (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[6] }), .b4_nUAi_0(
        b4_nUAi_288), .b4_nUAi_30(b4_nUAi_318), .b4_nUAi_27(
        b4_nUAi_315), .b4_nUAi_24(b4_nUAi_312), .b4_nUAi_21(
        b4_nUAi_309), .b4_nUAi_18(b4_nUAi_306), .b6_2ZTGIf_6(
        b6_2ZTGIf_102), .b6_2ZTGIf_4(b6_2ZTGIf_100), .b6_2ZTGIf_3(
        b6_2ZTGIf_99), .b6_2ZTGIf_2(b6_2ZTGIf_98), .b6_2ZTGIf_1(
        b6_2ZTGIf_97), .b6_2ZTGIf_0(b6_2ZTGIf_96), .b6_2ZTGIf_10(
        b6_2ZTGIf_106), .b6_2ZTGIf_9(b6_2ZTGIf_105), .b6_2ZTGIf_8(
        b6_2ZTGIf_104), .b6_2ZTGIf_7(b6_2ZTGIf_103), .N_25(N_25_35), 
        .N_27(N_27_35), .N_25_0(N_25_36), .N_27_0(N_27_36), .N_25_1(
        N_25_37), .N_27_1(N_27_37), .N_25_2(N_25_38), .N_27_2(N_27_38), 
        .N_25_3(N_25_39), .N_27_3(N_27_39), .N_25_4(N_25_40), .N_27_4(
        N_27_40));
    VCC VCC (.Y(VCC_net_1));
    b9_O2yyf_fG2_x_12_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_06 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[20] }), .b4_nUAi_0(
        b4_nUAi_960), .b4_nUAi_30(b4_nUAi_990), .b4_nUAi_27(
        b4_nUAi_987), .b4_nUAi_24(b4_nUAi_984), .b4_nUAi_21(
        b4_nUAi_981), .b4_nUAi_18(b4_nUAi_978), .b6_2ZTGIf_6(
        b6_2ZTGIf_326), .b6_2ZTGIf_4(b6_2ZTGIf_324), .b6_2ZTGIf_3(
        b6_2ZTGIf_323), .b6_2ZTGIf_2(b6_2ZTGIf_322), .b6_2ZTGIf_1(
        b6_2ZTGIf_321), .b6_2ZTGIf_0(b6_2ZTGIf_320), .b6_2ZTGIf_10(
        b6_2ZTGIf_330), .b6_2ZTGIf_9(b6_2ZTGIf_329), .b6_2ZTGIf_8(
        b6_2ZTGIf_328), .b6_2ZTGIf_7(b6_2ZTGIf_327), .N_25(N_25_119), 
        .N_27(N_27_119), .N_25_0(N_25_120), .N_27_0(N_27_120), .N_25_1(
        N_25_121), .N_27_1(N_27_121), .N_25_2(N_25_122), .N_27_2(
        N_27_122), .N_25_3(N_25_123), .N_27_3(N_27_123), .N_25_4(
        N_25_124), .N_27_4(N_27_124));
    SLE \b14_CZS0wfY_d_FH9m[0]  (.D(\b13_CZS0wfY_d_FH9[0] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[0]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[2]  (.D(\b13_CZS0wfY_d_FH9[2] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[2]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[20]  (.D(\b13_CZS0wfY_d_FH9[20] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[20]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[18]  (.D(\b13_CZS0wfY_d_FH9[18] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[18]_net_1 ));
    b9_O2yyf_fG2_x_9_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_0F (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[23] }), .b4_nUAi_18(
        b4_nUAi_1107), .b4_nUAi_12(b4_nUAi_1101), .b4_nUAi_6(
        b4_nUAi_1095), .b4_nUAi_0(b4_nUAi_1089), .b6_2ZTGIf_6(
        b6_2ZTGIf_375), .b6_2ZTGIf_4(b6_2ZTGIf_373), .b6_2ZTGIf_2(
        b6_2ZTGIf_371), .b6_2ZTGIf_0(b6_2ZTGIf_369), .N_25(N_25_137), 
        .N_27(N_27_137), .N_25_0(N_25_138), .N_27_0(N_27_138), .N_25_1(
        N_25_139), .N_27_1(N_27_139), .N_25_2(N_25_140), .N_27_2(
        N_27_140), .N_25_3(N_25_141), .b7_PSyi3wy(b7_PSyi3wy), .N_27_3(
        N_27_141));
    SLE \b14_CZS0wfY_d_FH9m[11]  (.D(\b13_CZS0wfY_d_FH9[11] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[11]_net_1 ));
    b9_O2yyf_fG2_x_16_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_aP (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[16] }), .b4_nUAi_0(
        b4_nUAi_768), .b4_nUAi_30(b4_nUAi_798), .b4_nUAi_27(
        b4_nUAi_795), .b4_nUAi_24(b4_nUAi_792), .b4_nUAi_21(
        b4_nUAi_789), .b4_nUAi_18(b4_nUAi_786), .b6_2ZTGIf_6(
        b6_2ZTGIf_262), .b6_2ZTGIf_4(b6_2ZTGIf_260), .b6_2ZTGIf_3(
        b6_2ZTGIf_259), .b6_2ZTGIf_2(b6_2ZTGIf_258), .b6_2ZTGIf_1(
        b6_2ZTGIf_257), .b6_2ZTGIf_0(b6_2ZTGIf_256), .b6_2ZTGIf_10(
        b6_2ZTGIf_266), .b6_2ZTGIf_9(b6_2ZTGIf_265), .b6_2ZTGIf_8(
        b6_2ZTGIf_264), .b6_2ZTGIf_7(b6_2ZTGIf_263), .N_25(N_25_95), 
        .N_27(N_27_95), .N_25_0(N_25_96), .N_27_0(N_27_96), .N_25_1(
        N_25_97), .N_27_1(N_27_97), .N_25_2(N_25_98), .N_27_2(N_27_98), 
        .N_25_3(N_25_99), .N_27_3(N_27_99), .N_25_4(N_25_100), .N_27_4(
        N_27_100));
    SLE \b14_CZS0wfY_d_FH9m[9]  (.D(\b13_CZS0wfY_d_FH9[9] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[9]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[22]  (.D(\b13_CZS0wfY_d_FH9[22] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[22]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[14]  (.D(\b13_CZS0wfY_d_FH9[14] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[14]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \b14_CZS0wfY_d_FH9m[16]  (.D(\b13_CZS0wfY_d_FH9[16] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[16]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[4]  (.D(\b13_CZS0wfY_d_FH9[4] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[4]_net_1 ));
    b9_O2yyf_fG2_x_20_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_aX (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[12] }), .b4_nUAi_0(
        b4_nUAi_576), .b4_nUAi_30(b4_nUAi_606), .b4_nUAi_27(
        b4_nUAi_603), .b4_nUAi_24(b4_nUAi_600), .b4_nUAi_21(
        b4_nUAi_597), .b4_nUAi_18(b4_nUAi_594), .b6_2ZTGIf_6(
        b6_2ZTGIf_198), .b6_2ZTGIf_4(b6_2ZTGIf_196), .b6_2ZTGIf_3(
        b6_2ZTGIf_195), .b6_2ZTGIf_2(b6_2ZTGIf_194), .b6_2ZTGIf_1(
        b6_2ZTGIf_193), .b6_2ZTGIf_0(b6_2ZTGIf_192), .b6_2ZTGIf_10(
        b6_2ZTGIf_202), .b6_2ZTGIf_9(b6_2ZTGIf_201), .b6_2ZTGIf_8(
        b6_2ZTGIf_200), .b6_2ZTGIf_7(b6_2ZTGIf_199), .N_25(N_25_71), 
        .N_27(N_27_71), .N_25_0(N_25_72), .N_27_0(N_27_72), .N_25_1(
        N_25_73), .N_27_1(N_27_73), .N_25_2(N_25_74), .N_27_2(N_27_74), 
        .N_25_3(N_25_75), .N_27_3(N_27_75), .N_25_4(N_25_76), .N_27_4(
        N_27_76));
    b9_O2yyf_fG2_x_21_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_a7 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[11] }), .b4_nUAi_0(
        b4_nUAi_528), .b4_nUAi_30(b4_nUAi_558), .b4_nUAi_27(
        b4_nUAi_555), .b4_nUAi_24(b4_nUAi_552), .b4_nUAi_21(
        b4_nUAi_549), .b4_nUAi_18(b4_nUAi_546), .b6_2ZTGIf_6(
        b6_2ZTGIf_182), .b6_2ZTGIf_4(b6_2ZTGIf_180), .b6_2ZTGIf_3(
        b6_2ZTGIf_179), .b6_2ZTGIf_2(b6_2ZTGIf_178), .b6_2ZTGIf_1(
        b6_2ZTGIf_177), .b6_2ZTGIf_0(b6_2ZTGIf_176), .b6_2ZTGIf_10(
        b6_2ZTGIf_186), .b6_2ZTGIf_9(b6_2ZTGIf_185), .b6_2ZTGIf_8(
        b6_2ZTGIf_184), .b6_2ZTGIf_7(b6_2ZTGIf_183), .N_25(N_25_65), 
        .N_27(N_27_65), .N_25_0(N_25_66), .N_27_0(N_27_66), .N_25_1(
        N_25_67), .N_27_1(N_27_67), .N_25_2(N_25_68), .N_27_2(N_27_68), 
        .N_25_3(N_25_69), .N_27_3(N_27_69), .N_25_4(N_25_70), .N_27_4(
        N_27_70));
    b9_O2yyf_fG2_x_32_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_9 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[0] }), .b4_nUAi_0(
        b4_nUAi_0), .b4_nUAi_30(b4_nUAi_30), .b4_nUAi_27(b4_nUAi_27), 
        .b4_nUAi_24(b4_nUAi_24), .b4_nUAi_21(b4_nUAi_21), .b4_nUAi_18(
        b4_nUAi_18), .b6_2ZTGIf_6(b6_2ZTGIf_6), .b6_2ZTGIf_4(
        b6_2ZTGIf_4), .b6_2ZTGIf_3(b6_2ZTGIf_3), .b6_2ZTGIf_2(
        b6_2ZTGIf_2), .b6_2ZTGIf_1(b6_2ZTGIf_1), .b6_2ZTGIf_0(
        b6_2ZTGIf_0), .b6_2ZTGIf_10(b6_2ZTGIf_10), .b6_2ZTGIf_9(
        b6_2ZTGIf_9), .b6_2ZTGIf_8(b6_2ZTGIf_8), .b6_2ZTGIf_7(
        b6_2ZTGIf_7), .N_25(N_25), .N_27(N_27), .N_25_0(N_25_0), 
        .N_27_0(N_27_0), .N_25_1(N_25_1), .N_27_1(N_27_1), .N_25_2(
        N_25_2), .N_27_2(N_27_2), .N_25_3(N_25_3), .N_27_3(N_27_3), 
        .N_25_4(N_25_4), .N_27_4(N_27_4));
    b9_O2yyf_fG2_x_31_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_a (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[1] }), .b4_nUAi_0(
        b4_nUAi_48), .b4_nUAi_30(b4_nUAi_78), .b4_nUAi_27(b4_nUAi_75), 
        .b4_nUAi_24(b4_nUAi_72), .b4_nUAi_21(b4_nUAi_69), .b4_nUAi_18(
        b4_nUAi_66), .b6_2ZTGIf_6(b6_2ZTGIf_22), .b6_2ZTGIf_4(
        b6_2ZTGIf_20), .b6_2ZTGIf_3(b6_2ZTGIf_19), .b6_2ZTGIf_2(
        b6_2ZTGIf_18), .b6_2ZTGIf_1(b6_2ZTGIf_17), .b6_2ZTGIf_0(
        b6_2ZTGIf_16), .b6_2ZTGIf_10(b6_2ZTGIf_26), .b6_2ZTGIf_9(
        b6_2ZTGIf_25), .b6_2ZTGIf_8(b6_2ZTGIf_24), .b6_2ZTGIf_7(
        b6_2ZTGIf_23), .N_25(N_25_5), .N_27(N_27_5), .N_25_0(N_25_6), 
        .N_27_0(N_27_6), .N_25_1(N_25_7), .N_27_1(N_27_7), .N_25_2(
        N_25_8), .N_27_2(N_27_8), .N_25_3(N_25_9), .N_27_3(N_27_9), 
        .N_25_4(N_25_10), .N_27_4(N_27_10));
    b9_O2yyf_fG2_x_0_0 b25_O2yyf_fG2_MiQA1E6_p_lnxob (
        .b14_CZS0wfY_d_FH9m({\b14_CZS0wfY_d_FH9m[23]_net_1 , 
        \b14_CZS0wfY_d_FH9m[22]_net_1 , \b14_CZS0wfY_d_FH9m[21]_net_1 , 
        \b14_CZS0wfY_d_FH9m[20]_net_1 , \b14_CZS0wfY_d_FH9m[19]_net_1 , 
        \b14_CZS0wfY_d_FH9m[18]_net_1 , \b14_CZS0wfY_d_FH9m[17]_net_1 , 
        \b14_CZS0wfY_d_FH9m[16]_net_1 , \b14_CZS0wfY_d_FH9m[15]_net_1 , 
        \b14_CZS0wfY_d_FH9m[14]_net_1 , \b14_CZS0wfY_d_FH9m[13]_net_1 , 
        \b14_CZS0wfY_d_FH9m[12]_net_1 , \b14_CZS0wfY_d_FH9m[11]_net_1 , 
        \b14_CZS0wfY_d_FH9m[10]_net_1 , \b14_CZS0wfY_d_FH9m[9]_net_1 , 
        \b14_CZS0wfY_d_FH9m[8]_net_1 , \b14_CZS0wfY_d_FH9m[7]_net_1 , 
        \b14_CZS0wfY_d_FH9m[6]_net_1 , \b14_CZS0wfY_d_FH9m[5]_net_1 , 
        \b14_CZS0wfY_d_FH9m[4]_net_1 , \b14_CZS0wfY_d_FH9m[3]_net_1 , 
        \b14_CZS0wfY_d_FH9m[2]_net_1 , \b14_CZS0wfY_d_FH9m[1]_net_1 , 
        \b14_CZS0wfY_d_FH9m[0]_net_1 }), .b11_uUT0JC4gFrY({
        b11_uUT0JC4gFrY[1]}));
    SLE \b14_CZS0wfY_d_FH9m[21]  (.D(\b13_CZS0wfY_d_FH9[21] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[21]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[8]  (.D(\b13_CZS0wfY_d_FH9[8] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[8]_net_1 ));
    b9_O2yyf_fG2_x_27_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_c (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[5] }), .b4_nUAi_0(
        b4_nUAi_240), .b4_nUAi_30(b4_nUAi_270), .b4_nUAi_27(
        b4_nUAi_267), .b4_nUAi_24(b4_nUAi_264), .b4_nUAi_21(
        b4_nUAi_261), .b4_nUAi_18(b4_nUAi_258), .b6_2ZTGIf_6(
        b6_2ZTGIf_86), .b6_2ZTGIf_4(b6_2ZTGIf_84), .b6_2ZTGIf_3(
        b6_2ZTGIf_83), .b6_2ZTGIf_2(b6_2ZTGIf_82), .b6_2ZTGIf_1(
        b6_2ZTGIf_81), .b6_2ZTGIf_0(b6_2ZTGIf_80), .b6_2ZTGIf_10(
        b6_2ZTGIf_90), .b6_2ZTGIf_9(b6_2ZTGIf_89), .b6_2ZTGIf_8(
        b6_2ZTGIf_88), .b6_2ZTGIf_7(b6_2ZTGIf_87), .N_25(N_25_29), 
        .N_27(N_27_29), .N_25_0(N_25_30), .N_27_0(N_27_30), .N_25_1(
        N_25_31), .N_27_1(N_27_31), .N_25_2(N_25_32), .N_27_2(N_27_32), 
        .N_25_3(N_25_33), .N_27_3(N_27_33), .N_25_4(N_25_34), .N_27_4(
        N_27_34));
    b9_O2yyf_fG2_x_28_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_8 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[4] }), .b4_nUAi_0(
        b4_nUAi_192), .b4_nUAi_30(b4_nUAi_222), .b4_nUAi_27(
        b4_nUAi_219), .b4_nUAi_24(b4_nUAi_216), .b4_nUAi_21(
        b4_nUAi_213), .b4_nUAi_18(b4_nUAi_210), .b6_2ZTGIf_6(
        b6_2ZTGIf_70), .b6_2ZTGIf_4(b6_2ZTGIf_68), .b6_2ZTGIf_3(
        b6_2ZTGIf_67), .b6_2ZTGIf_2(b6_2ZTGIf_66), .b6_2ZTGIf_1(
        b6_2ZTGIf_65), .b6_2ZTGIf_0(b6_2ZTGIf_64), .b6_2ZTGIf_10(
        b6_2ZTGIf_74), .b6_2ZTGIf_9(b6_2ZTGIf_73), .b6_2ZTGIf_8(
        b6_2ZTGIf_72), .b6_2ZTGIf_7(b6_2ZTGIf_71), .N_25(N_25_23), 
        .N_27(N_27_23), .N_25_0(N_25_24), .N_27_0(N_27_24), .N_25_1(
        N_25_25), .N_27_1(N_27_25), .N_25_2(N_25_26), .N_27_2(N_27_26), 
        .N_25_3(N_25_27), .N_27_3(N_27_27), .N_25_4(N_25_28), .N_27_4(
        N_27_28));
    b9_O2yyf_fG2_x_10_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_0X (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[22] }), .b4_nUAi_0(
        b4_nUAi_1056), .b4_nUAi_30(b4_nUAi_1086), .b4_nUAi_27(
        b4_nUAi_1083), .b4_nUAi_24(b4_nUAi_1080), .b4_nUAi_21(
        b4_nUAi_1077), .b4_nUAi_18(b4_nUAi_1074), .b6_2ZTGIf_6(
        b6_2ZTGIf_358), .b6_2ZTGIf_4(b6_2ZTGIf_356), .b6_2ZTGIf_3(
        b6_2ZTGIf_355), .b6_2ZTGIf_2(b6_2ZTGIf_354), .b6_2ZTGIf_1(
        b6_2ZTGIf_353), .b6_2ZTGIf_0(b6_2ZTGIf_352), .b6_2ZTGIf_10(
        b6_2ZTGIf_362), .b6_2ZTGIf_9(b6_2ZTGIf_361), .b6_2ZTGIf_8(
        b6_2ZTGIf_360), .b6_2ZTGIf_7(b6_2ZTGIf_359), .N_25(N_25_131), 
        .N_27(N_27_131), .N_25_0(N_25_132), .N_27_0(N_27_132), .N_25_1(
        N_25_133), .N_27_1(N_27_133), .N_25_2(N_25_134), .N_27_2(
        N_27_134), .N_25_3(N_25_135), .N_27_3(N_27_135), .N_25_4(
        N_25_136), .N_27_4(N_27_136));
    b9_O2yyf_fG2_x_11_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_07 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[21] }), .b4_nUAi_0(
        b4_nUAi_1008), .b4_nUAi_30(b4_nUAi_1038), .b4_nUAi_27(
        b4_nUAi_1035), .b4_nUAi_24(b4_nUAi_1032), .b4_nUAi_21(
        b4_nUAi_1029), .b4_nUAi_18(b4_nUAi_1026), .b6_2ZTGIf_6(
        b6_2ZTGIf_342), .b6_2ZTGIf_4(b6_2ZTGIf_340), .b6_2ZTGIf_3(
        b6_2ZTGIf_339), .b6_2ZTGIf_2(b6_2ZTGIf_338), .b6_2ZTGIf_1(
        b6_2ZTGIf_337), .b6_2ZTGIf_0(b6_2ZTGIf_336), .b6_2ZTGIf_10(
        b6_2ZTGIf_346), .b6_2ZTGIf_9(b6_2ZTGIf_345), .b6_2ZTGIf_8(
        b6_2ZTGIf_344), .b6_2ZTGIf_7(b6_2ZTGIf_343), .N_25(N_25_125), 
        .N_27(N_27_125), .N_25_0(N_25_126), .N_27_0(N_27_126), .N_25_1(
        N_25_127), .N_27_1(N_27_127), .N_25_2(N_25_128), .N_27_2(
        N_27_128), .N_25_3(N_25_129), .N_27_3(N_27_129), .N_25_4(
        N_25_130), .N_27_4(N_27_130));
    b9_O2yyf_fG2_x_24_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_F (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[8] }), .b4_nUAi_0(
        b4_nUAi_384), .b4_nUAi_30(b4_nUAi_414), .b4_nUAi_27(
        b4_nUAi_411), .b4_nUAi_24(b4_nUAi_408), .b4_nUAi_21(
        b4_nUAi_405), .b4_nUAi_18(b4_nUAi_402), .b6_2ZTGIf_6(
        b6_2ZTGIf_134), .b6_2ZTGIf_4(b6_2ZTGIf_132), .b6_2ZTGIf_3(
        b6_2ZTGIf_131), .b6_2ZTGIf_2(b6_2ZTGIf_130), .b6_2ZTGIf_1(
        b6_2ZTGIf_129), .b6_2ZTGIf_0(b6_2ZTGIf_128), .b6_2ZTGIf_10(
        b6_2ZTGIf_138), .b6_2ZTGIf_9(b6_2ZTGIf_137), .b6_2ZTGIf_8(
        b6_2ZTGIf_136), .b6_2ZTGIf_7(b6_2ZTGIf_135), .N_25(N_25_47), 
        .N_27(N_27_47), .N_25_0(N_25_48), .N_27_0(N_27_48), .N_25_1(
        N_25_49), .N_27_1(N_27_49), .N_25_2(N_25_50), .N_27_2(N_27_50), 
        .N_25_3(N_25_51), .N_27_3(N_27_51), .N_25_4(N_25_52), .N_27_4(
        N_27_52));
    b9_O2yyf_fG2_x_13_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_aa (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[19] }), .b4_nUAi_0(
        b4_nUAi_912), .b4_nUAi_30(b4_nUAi_942), .b4_nUAi_27(
        b4_nUAi_939), .b4_nUAi_24(b4_nUAi_936), .b4_nUAi_21(
        b4_nUAi_933), .b4_nUAi_18(b4_nUAi_930), .b6_2ZTGIf_6(
        b6_2ZTGIf_310), .b6_2ZTGIf_4(b6_2ZTGIf_308), .b6_2ZTGIf_3(
        b6_2ZTGIf_307), .b6_2ZTGIf_2(b6_2ZTGIf_306), .b6_2ZTGIf_1(
        b6_2ZTGIf_305), .b6_2ZTGIf_0(b6_2ZTGIf_304), .b6_2ZTGIf_10(
        b6_2ZTGIf_314), .b6_2ZTGIf_9(b6_2ZTGIf_313), .b6_2ZTGIf_8(
        b6_2ZTGIf_312), .b6_2ZTGIf_7(b6_2ZTGIf_311), .N_25(N_25_113), 
        .N_27(N_27_113), .N_25_0(N_25_114), .N_27_0(N_27_114), .N_25_1(
        N_25_115), .N_27_1(N_27_115), .N_25_2(N_25_116), .N_27_2(
        N_27_116), .N_25_3(N_25_117), .N_27_3(N_27_117), .N_25_4(
        N_25_118), .N_27_4(N_27_118));
    b9_O2yyf_fG2_x_15_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_aY (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[17] }), .b4_nUAi_0(
        b4_nUAi_816), .b4_nUAi_30(b4_nUAi_846), .b4_nUAi_27(
        b4_nUAi_843), .b4_nUAi_24(b4_nUAi_840), .b4_nUAi_21(
        b4_nUAi_837), .b4_nUAi_18(b4_nUAi_834), .b6_2ZTGIf_6(
        b6_2ZTGIf_278), .b6_2ZTGIf_4(b6_2ZTGIf_276), .b6_2ZTGIf_3(
        b6_2ZTGIf_275), .b6_2ZTGIf_2(b6_2ZTGIf_274), .b6_2ZTGIf_1(
        b6_2ZTGIf_273), .b6_2ZTGIf_0(b6_2ZTGIf_272), .b6_2ZTGIf_10(
        b6_2ZTGIf_282), .b6_2ZTGIf_9(b6_2ZTGIf_281), .b6_2ZTGIf_8(
        b6_2ZTGIf_280), .b6_2ZTGIf_7(b6_2ZTGIf_279), .N_25(N_25_101), 
        .N_27(N_27_101), .N_25_0(N_25_102), .N_27_0(N_27_102), .N_25_1(
        N_25_103), .N_27_1(N_27_103), .N_25_2(N_25_104), .N_27_2(
        N_27_104), .N_25_3(N_25_105), .N_27_3(N_27_105), .N_25_4(
        N_25_106), .N_27_4(N_27_106));
    SLE \b14_CZS0wfY_d_FH9m[5]  (.D(\b13_CZS0wfY_d_FH9[5] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[5]_net_1 ));
    b9_O2yyf_fG2_x_18_0 b28_O2yyf_fG2_MiQA1E6_r_lnxob_a5 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[14] }), .b4_nUAi_0(
        b4_nUAi_672), .b4_nUAi_30(b4_nUAi_702), .b4_nUAi_27(
        b4_nUAi_699), .b4_nUAi_24(b4_nUAi_696), .b4_nUAi_21(
        b4_nUAi_693), .b4_nUAi_18(b4_nUAi_690), .b6_2ZTGIf_6(
        b6_2ZTGIf_230), .b6_2ZTGIf_4(b6_2ZTGIf_228), .b6_2ZTGIf_3(
        b6_2ZTGIf_227), .b6_2ZTGIf_2(b6_2ZTGIf_226), .b6_2ZTGIf_1(
        b6_2ZTGIf_225), .b6_2ZTGIf_0(b6_2ZTGIf_224), .b6_2ZTGIf_10(
        b6_2ZTGIf_234), .b6_2ZTGIf_9(b6_2ZTGIf_233), .b6_2ZTGIf_8(
        b6_2ZTGIf_232), .b6_2ZTGIf_7(b6_2ZTGIf_231), .N_25(N_25_83), 
        .N_27(N_27_83), .N_25_0(N_25_84), .N_27_0(N_27_84), .N_25_1(
        N_25_85), .N_27_1(N_27_85), .N_25_2(N_25_86), .N_27_2(N_27_86), 
        .N_25_3(N_25_87), .N_27_3(N_27_87), .N_25_4(N_25_88), .N_27_4(
        N_27_88));
    b9_O2yyf_fG2_x_30_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_0 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[2] }), .b4_nUAi_0(
        b4_nUAi_96), .b4_nUAi_30(b4_nUAi_126), .b4_nUAi_27(b4_nUAi_123)
        , .b4_nUAi_24(b4_nUAi_120), .b4_nUAi_21(b4_nUAi_117), 
        .b4_nUAi_18(b4_nUAi_114), .b6_2ZTGIf_6(b6_2ZTGIf_38), 
        .b6_2ZTGIf_4(b6_2ZTGIf_36), .b6_2ZTGIf_3(b6_2ZTGIf_35), 
        .b6_2ZTGIf_2(b6_2ZTGIf_34), .b6_2ZTGIf_1(b6_2ZTGIf_33), 
        .b6_2ZTGIf_0(b6_2ZTGIf_32), .b6_2ZTGIf_10(b6_2ZTGIf_42), 
        .b6_2ZTGIf_9(b6_2ZTGIf_41), .b6_2ZTGIf_8(b6_2ZTGIf_40), 
        .b6_2ZTGIf_7(b6_2ZTGIf_39), .N_25(N_25_11), .N_27(N_27_11), 
        .N_25_0(N_25_12), .N_27_0(N_27_12), .N_25_1(N_25_13), .N_27_1(
        N_27_13), .N_25_2(N_25_14), .N_27_2(N_27_14), .N_25_3(N_25_15), 
        .N_27_3(N_27_15), .N_25_4(N_25_16), .N_27_4(N_27_16));
    SLE \b14_CZS0wfY_d_FH9m[13]  (.D(\b13_CZS0wfY_d_FH9[13] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[13]_net_1 ));
    b9_O2yyf_fG2_x_25_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_1 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[7] }), .b4_nUAi_0(
        b4_nUAi_336), .b4_nUAi_30(b4_nUAi_366), .b4_nUAi_27(
        b4_nUAi_363), .b4_nUAi_24(b4_nUAi_360), .b4_nUAi_21(
        b4_nUAi_357), .b4_nUAi_18(b4_nUAi_354), .b6_2ZTGIf_6(
        b6_2ZTGIf_118), .b6_2ZTGIf_4(b6_2ZTGIf_116), .b6_2ZTGIf_3(
        b6_2ZTGIf_115), .b6_2ZTGIf_2(b6_2ZTGIf_114), .b6_2ZTGIf_1(
        b6_2ZTGIf_113), .b6_2ZTGIf_0(b6_2ZTGIf_112), .b6_2ZTGIf_10(
        b6_2ZTGIf_122), .b6_2ZTGIf_9(b6_2ZTGIf_121), .b6_2ZTGIf_8(
        b6_2ZTGIf_120), .b6_2ZTGIf_7(b6_2ZTGIf_119), .N_25(N_25_41), 
        .N_27(N_27_41), .N_25_0(N_25_42), .N_27_0(N_27_42), .N_25_1(
        N_25_43), .N_27_1(N_27_43), .N_25_2(N_25_44), .N_27_2(N_27_44), 
        .N_25_3(N_25_45), .N_27_3(N_27_45), .N_25_4(N_25_46), .N_27_4(
        N_27_46));
    SLE \b14_CZS0wfY_d_FH9m[6]  (.D(\b13_CZS0wfY_d_FH9[6] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[6]_net_1 ));
    b9_O2yyf_fG2_x_23_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_d (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[9] }), .b4_nUAi_0(
        b4_nUAi_432), .b4_nUAi_30(b4_nUAi_462), .b4_nUAi_27(
        b4_nUAi_459), .b4_nUAi_24(b4_nUAi_456), .b4_nUAi_21(
        b4_nUAi_453), .b4_nUAi_18(b4_nUAi_450), .b6_2ZTGIf_6(
        b6_2ZTGIf_150), .b6_2ZTGIf_4(b6_2ZTGIf_148), .b6_2ZTGIf_3(
        b6_2ZTGIf_147), .b6_2ZTGIf_2(b6_2ZTGIf_146), .b6_2ZTGIf_1(
        b6_2ZTGIf_145), .b6_2ZTGIf_0(b6_2ZTGIf_144), .b6_2ZTGIf_10(
        b6_2ZTGIf_154), .b6_2ZTGIf_9(b6_2ZTGIf_153), .b6_2ZTGIf_8(
        b6_2ZTGIf_152), .b6_2ZTGIf_7(b6_2ZTGIf_151), .N_25(N_25_53), 
        .N_27(N_27_53), .N_25_0(N_25_54), .N_27_0(N_27_54), .N_25_1(
        N_25_55), .N_27_1(N_27_55), .N_25_2(N_25_56), .N_27_2(N_27_56), 
        .N_25_3(N_25_57), .N_27_3(N_27_57), .N_25_4(N_25_58), .N_27_4(
        N_27_58));
    SLE \b14_CZS0wfY_d_FH9m[1]  (.D(\b13_CZS0wfY_d_FH9[1] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[1]_net_1 ));
    
endmodule


module b8_1LbcQDr1_x_51_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [325:325] mdiclink_reg;
input  [51:51] b11_OFWNT9L_8tZ;
input  [976:975] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[325]), .B(
        b11_OFWNT9L_8tZ[51]), .C(b4_nUAi[976]), .D(b4_nUAi[975]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[325]), .B(
        b11_OFWNT9L_8tZ[51]), .C(b4_nUAi[976]), .D(b4_nUAi[975]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_326_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [50:50] mdiclink_reg;
input  [326:326] b11_OFWNT9L_8tZ;
input  [152:150] b4_nUAi;
output [50:50] b6_2ZTGIf;

    wire b3_P_F_6_bm_190, b3_P_F_6_am_190, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_190), .B(
        b4_nUAi[152]), .C(b3_P_F_6_am_190), .Y(b6_2ZTGIf[50]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[50]), .B(
        b11_OFWNT9L_8tZ[326]), .C(b4_nUAi[151]), .D(b4_nUAi[150]), .Y(
        b3_P_F_6_am_190));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[50]), .B(
        b11_OFWNT9L_8tZ[326]), .C(b4_nUAi[150]), .D(b4_nUAi[151]), .Y(
        b3_P_F_6_bm_190));
    
endmodule


module b8_1LbcQDr1_x_294_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [82:82] mdiclink_reg;
input  [294:294] b11_OFWNT9L_8tZ;
input  [248:246] b4_nUAi;
output [82:82] b6_2ZTGIf;

    wire b3_P_F_6_bm_210, b3_P_F_6_am_210, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_210), .B(
        b4_nUAi[248]), .C(b3_P_F_6_am_210), .Y(b6_2ZTGIf[82]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[82]), .B(
        b11_OFWNT9L_8tZ[294]), .C(b4_nUAi[247]), .D(b4_nUAi[246]), .Y(
        b3_P_F_6_am_210));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[82]), .B(
        b11_OFWNT9L_8tZ[294]), .C(b4_nUAi[246]), .D(b4_nUAi[247]), .Y(
        b3_P_F_6_bm_210));
    
endmodule


module b8_1LbcQDr1_x_8_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [368:368] mdiclink_reg;
input  [8:8] b11_OFWNT9L_8tZ;
input  [1105:1104] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[368]), .B(
        b11_OFWNT9L_8tZ[8]), .C(b4_nUAi[1105]), .D(b4_nUAi[1104]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[368]), .B(
        b11_OFWNT9L_8tZ[8]), .C(b4_nUAi[1105]), .D(b4_nUAi[1104]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_65_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [311:311] mdiclink_reg;
input  [65:65] b11_OFWNT9L_8tZ;
input  [935:933] b4_nUAi;
output [311:311] b6_2ZTGIf;

    wire b3_P_F_6_bm_112, b3_P_F_6_am_112, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_112), .B(
        b4_nUAi[935]), .C(b3_P_F_6_am_112), .Y(b6_2ZTGIf[311]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[311]), .B(
        b11_OFWNT9L_8tZ[65]), .C(b4_nUAi[934]), .D(b4_nUAi[933]), .Y(
        b3_P_F_6_am_112));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[311]), .B(
        b11_OFWNT9L_8tZ[65]), .C(b4_nUAi[933]), .D(b4_nUAi[934]), .Y(
        b3_P_F_6_bm_112));
    
endmodule


module b8_1LbcQDr1_x_75_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [301:301] mdiclink_reg;
input  [75:75] b11_OFWNT9L_8tZ;
input  [904:903] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[301]), .B(
        b11_OFWNT9L_8tZ[75]), .C(b4_nUAi[904]), .D(b4_nUAi[903]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[301]), .B(
        b11_OFWNT9L_8tZ[75]), .C(b4_nUAi[904]), .D(b4_nUAi[903]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_138_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [238:238] mdiclink_reg;
input  [138:138] b11_OFWNT9L_8tZ;
input  [715:714] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[238]), .B(
        b11_OFWNT9L_8tZ[138]), .C(b4_nUAi[715]), .D(b4_nUAi[714]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[238]), .B(
        b11_OFWNT9L_8tZ[138]), .C(b4_nUAi[715]), .D(b4_nUAi[714]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_255_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [121:121] mdiclink_reg;
input  [255:255] b11_OFWNT9L_8tZ;
input  [365:363] b4_nUAi;
output [121:121] b6_2ZTGIf;

    wire b3_P_F_6_bm_10, b3_P_F_6_am_10, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_10), .B(
        b4_nUAi[365]), .C(b3_P_F_6_am_10), .Y(b6_2ZTGIf[121]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[121]), .B(
        b11_OFWNT9L_8tZ[255]), .C(b4_nUAi[364]), .D(b4_nUAi[363]), .Y(
        b3_P_F_6_am_10));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[121]), .B(
        b11_OFWNT9L_8tZ[255]), .C(b4_nUAi[363]), .D(b4_nUAi[364]), .Y(
        b3_P_F_6_bm_10));
    
endmodule


module b8_1LbcQDr1_x_92_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [284:284] mdiclink_reg;
input  [92:92] b11_OFWNT9L_8tZ;
input  [853:852] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[284]), .B(
        b11_OFWNT9L_8tZ[92]), .C(b4_nUAi[853]), .D(b4_nUAi[852]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[284]), .B(
        b11_OFWNT9L_8tZ[92]), .C(b4_nUAi[853]), .D(b4_nUAi[852]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_28_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [348:348] mdiclink_reg;
input  [28:28] b11_OFWNT9L_8tZ;
input  [1045:1044] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[348]), .B(
        b11_OFWNT9L_8tZ[28]), .C(b4_nUAi[1045]), .D(b4_nUAi[1044]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[348]), .B(
        b11_OFWNT9L_8tZ[28]), .C(b4_nUAi[1045]), .D(b4_nUAi[1044]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_54_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [322:322] mdiclink_reg;
input  [54:54] b11_OFWNT9L_8tZ;
input  [968:966] b4_nUAi;
output [322:322] b6_2ZTGIf;

    wire b3_P_F_6_bm_126, b3_P_F_6_am_126, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_126), .B(
        b4_nUAi[968]), .C(b3_P_F_6_am_126), .Y(b6_2ZTGIf[322]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[322]), .B(
        b11_OFWNT9L_8tZ[54]), .C(b4_nUAi[967]), .D(b4_nUAi[966]), .Y(
        b3_P_F_6_am_126));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[322]), .B(
        b11_OFWNT9L_8tZ[54]), .C(b4_nUAi[966]), .D(b4_nUAi[967]), .Y(
        b3_P_F_6_bm_126));
    
endmodule


module b8_1LbcQDr1_x_201_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [175:175] mdiclink_reg;
input  [201:201] b11_OFWNT9L_8tZ;
input  [526:525] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[175]), .B(
        b11_OFWNT9L_8tZ[201]), .C(b4_nUAi[526]), .D(b4_nUAi[525]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[175]), .B(
        b11_OFWNT9L_8tZ[201]), .C(b4_nUAi[526]), .D(b4_nUAi[525]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_17_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [359:359] mdiclink_reg;
input  [17:17] b11_OFWNT9L_8tZ;
input  [1079:1077] b4_nUAi;
output [359:359] b6_2ZTGIf;

    wire b3_P_F_6_bm_142, b3_P_F_6_am_142, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_142), .B(
        b4_nUAi[1079]), .C(b3_P_F_6_am_142), .Y(b6_2ZTGIf[359]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[359]), .B(
        b11_OFWNT9L_8tZ[17]), .C(b4_nUAi[1078]), .D(b4_nUAi[1077]), .Y(
        b3_P_F_6_am_142));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[359]), .B(
        b11_OFWNT9L_8tZ[17]), .C(b4_nUAi[1077]), .D(b4_nUAi[1078]), .Y(
        b3_P_F_6_bm_142));
    
endmodule


module b8_1LbcQDr1_x_351_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [25:25] mdiclink_reg;
input  [351:351] b11_OFWNT9L_8tZ;
input  [77:75] b4_nUAi;
output [25:25] b6_2ZTGIf;

    wire b3_P_F_6_bm_164, b3_P_F_6_am_164, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_164), .B(
        b4_nUAi[77]), .C(b3_P_F_6_am_164), .Y(b6_2ZTGIf[25]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[25]), .B(
        b11_OFWNT9L_8tZ[351]), .C(b4_nUAi[76]), .D(b4_nUAi[75]), .Y(
        b3_P_F_6_am_164));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[25]), .B(
        b11_OFWNT9L_8tZ[351]), .C(b4_nUAi[75]), .D(b4_nUAi[76]), .Y(
        b3_P_F_6_bm_164));
    
endmodule


module b8_1LbcQDr1_x_311_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [65:65] mdiclink_reg;
input  [311:311] b11_OFWNT9L_8tZ;
input  [197:195] b4_nUAi;
output [65:65] b6_2ZTGIf;

    wire b3_P_F_6_bm_201, b3_P_F_6_am_201, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_201), .B(
        b4_nUAi[197]), .C(b3_P_F_6_am_201), .Y(b6_2ZTGIf[65]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[65]), .B(
        b11_OFWNT9L_8tZ[311]), .C(b4_nUAi[196]), .D(b4_nUAi[195]), .Y(
        b3_P_F_6_am_201));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[65]), .B(
        b11_OFWNT9L_8tZ[311]), .C(b4_nUAi[195]), .D(b4_nUAi[196]), .Y(
        b3_P_F_6_bm_201));
    
endmodule


module b8_1LbcQDr1_x_163_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [213:213] mdiclink_reg;
input  [163:163] b11_OFWNT9L_8tZ;
input  [640:639] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[213]), .B(
        b11_OFWNT9L_8tZ[163]), .C(b4_nUAi[640]), .D(b4_nUAi[639]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[213]), .B(
        b11_OFWNT9L_8tZ[163]), .C(b4_nUAi[640]), .D(b4_nUAi[639]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_342_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [34:34] mdiclink_reg;
input  [342:342] b11_OFWNT9L_8tZ;
input  [104:102] b4_nUAi;
output [34:34] b6_2ZTGIf;

    wire b3_P_F_6_bm_180, b3_P_F_6_am_180, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_180), .B(
        b4_nUAi[104]), .C(b3_P_F_6_am_180), .Y(b6_2ZTGIf[34]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[34]), .B(
        b11_OFWNT9L_8tZ[342]), .C(b4_nUAi[103]), .D(b4_nUAi[102]), .Y(
        b3_P_F_6_am_180));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[34]), .B(
        b11_OFWNT9L_8tZ[342]), .C(b4_nUAi[102]), .D(b4_nUAi[103]), .Y(
        b3_P_F_6_bm_180));
    
endmodule


module b8_1LbcQDr1_x_212_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [164:164] mdiclink_reg;
input  [212:212] b11_OFWNT9L_8tZ;
input  [494:492] b4_nUAi;
output [164:164] b6_2ZTGIf;

    wire b3_P_F_6_bm_44, b3_P_F_6_am_44, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_44), .B(
        b4_nUAi[494]), .C(b3_P_F_6_am_44), .Y(b6_2ZTGIf[164]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[164]), .B(
        b11_OFWNT9L_8tZ[212]), .C(b4_nUAi[493]), .D(b4_nUAi[492]), .Y(
        b3_P_F_6_am_44));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[164]), .B(
        b11_OFWNT9L_8tZ[212]), .C(b4_nUAi[492]), .D(b4_nUAi[493]), .Y(
        b3_P_F_6_bm_44));
    
endmodule


module b8_1LbcQDr1_x_42_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [334:334] mdiclink_reg;
input  [42:42] b11_OFWNT9L_8tZ;
input  [1003:1002] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[334]), .B(
        b11_OFWNT9L_8tZ[42]), .C(b4_nUAi[1003]), .D(b4_nUAi[1002]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[334]), .B(
        b11_OFWNT9L_8tZ[42]), .C(b4_nUAi[1003]), .D(b4_nUAi[1002]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_173_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [203:203] mdiclink_reg;
input  [173:173] b11_OFWNT9L_8tZ;
input  [610:609] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[203]), .B(
        b11_OFWNT9L_8tZ[173]), .C(b4_nUAi[610]), .D(b4_nUAi[609]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[203]), .B(
        b11_OFWNT9L_8tZ[173]), .C(b4_nUAi[610]), .D(b4_nUAi[609]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_210_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [166:166] mdiclink_reg;
input  [210:210] b11_OFWNT9L_8tZ;
input  [500:498] b4_nUAi;
output [166:166] b6_2ZTGIf;

    wire b3_P_F_6_bm_43, b3_P_F_6_am_43, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_43), .B(
        b4_nUAi[500]), .C(b3_P_F_6_am_43), .Y(b6_2ZTGIf[166]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[166]), .B(
        b11_OFWNT9L_8tZ[210]), .C(b4_nUAi[499]), .D(b4_nUAi[498]), .Y(
        b3_P_F_6_am_43));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[166]), .B(
        b11_OFWNT9L_8tZ[210]), .C(b4_nUAi[498]), .D(b4_nUAi[499]), .Y(
        b3_P_F_6_bm_43));
    
endmodule


module b8_1LbcQDr1_x_312_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [64:64] mdiclink_reg;
input  [312:312] b11_OFWNT9L_8tZ;
input  [194:192] b4_nUAi;
output [64:64] b6_2ZTGIf;

    wire b3_P_F_6_bm_202, b3_P_F_6_am_202, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_202), .B(
        b4_nUAi[194]), .C(b3_P_F_6_am_202), .Y(b6_2ZTGIf[64]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[64]), .B(
        b11_OFWNT9L_8tZ[312]), .C(b4_nUAi[193]), .D(b4_nUAi[192]), .Y(
        b3_P_F_6_am_202));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[64]), .B(
        b11_OFWNT9L_8tZ[312]), .C(b4_nUAi[192]), .D(b4_nUAi[193]), .Y(
        b3_P_F_6_bm_202));
    
endmodule


module b8_1LbcQDr1_x_82_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [294:294] mdiclink_reg;
input  [82:82] b11_OFWNT9L_8tZ;
input  [884:882] b4_nUAi;
output [294:294] b6_2ZTGIf;

    wire b3_P_F_6_bm_103, b3_P_F_6_am_103, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_103), .B(
        b4_nUAi[884]), .C(b3_P_F_6_am_103), .Y(b6_2ZTGIf[294]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[294]), .B(
        b11_OFWNT9L_8tZ[82]), .C(b4_nUAi[883]), .D(b4_nUAi[882]), .Y(
        b3_P_F_6_am_103));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[294]), .B(
        b11_OFWNT9L_8tZ[82]), .C(b4_nUAi[882]), .D(b4_nUAi[883]), .Y(
        b3_P_F_6_bm_103));
    
endmodule


module b8_1LbcQDr1_x_146_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [230:230] mdiclink_reg;
input  [146:146] b11_OFWNT9L_8tZ;
input  [692:690] b4_nUAi;
output [230:230] b6_2ZTGIf;

    wire b3_P_F_6_bm_217, b3_P_F_6_am_217, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_217), .B(
        b4_nUAi[692]), .C(b3_P_F_6_am_217), .Y(b6_2ZTGIf[230]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[230]), .B(
        b11_OFWNT9L_8tZ[146]), .C(b4_nUAi[691]), .D(b4_nUAi[690]), .Y(
        b3_P_F_6_am_217));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[230]), .B(
        b11_OFWNT9L_8tZ[146]), .C(b4_nUAi[690]), .D(b4_nUAi[691]), .Y(
        b3_P_F_6_bm_217));
    
endmodule


module b8_1LbcQDr1_x_197_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [179:179] mdiclink_reg;
input  [197:197] b11_OFWNT9L_8tZ;
input  [539:537] b4_nUAi;
output [179:179] b6_2ZTGIf;

    wire b3_P_F_6_bm_55, b3_P_F_6_am_55, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_55), .B(
        b4_nUAi[539]), .C(b3_P_F_6_am_55), .Y(b6_2ZTGIf[179]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[179]), .B(
        b11_OFWNT9L_8tZ[197]), .C(b4_nUAi[538]), .D(b4_nUAi[537]), .Y(
        b3_P_F_6_am_55));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[179]), .B(
        b11_OFWNT9L_8tZ[197]), .C(b4_nUAi[537]), .D(b4_nUAi[538]), .Y(
        b3_P_F_6_bm_55));
    
endmodule


module b8_1LbcQDr1_x_125_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [251:251] mdiclink_reg;
input  [125:125] b11_OFWNT9L_8tZ;
input  [754:753] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[251]), .B(
        b11_OFWNT9L_8tZ[125]), .C(b4_nUAi[754]), .D(b4_nUAi[753]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[251]), .B(
        b11_OFWNT9L_8tZ[125]), .C(b4_nUAi[754]), .D(b4_nUAi[753]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_232_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [144:144] mdiclink_reg;
input  [232:232] b11_OFWNT9L_8tZ;
input  [434:432] b4_nUAi;
output [144:144] b6_2ZTGIf;

    wire b3_P_F_6_bm_38, b3_P_F_6_am_38, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_38), .B(
        b4_nUAi[434]), .C(b3_P_F_6_am_38), .Y(b6_2ZTGIf[144]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[144]), .B(
        b11_OFWNT9L_8tZ[232]), .C(b4_nUAi[433]), .D(b4_nUAi[432]), .Y(
        b3_P_F_6_am_38));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[144]), .B(
        b11_OFWNT9L_8tZ[232]), .C(b4_nUAi[432]), .D(b4_nUAi[433]), .Y(
        b3_P_F_6_bm_38));
    
endmodule


module b8_1LbcQDr1_x_46_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [330:330] mdiclink_reg;
input  [46:46] b11_OFWNT9L_8tZ;
input  [992:990] b4_nUAi;
output [330:330] b6_2ZTGIf;

    wire b3_P_F_6_bm_119, b3_P_F_6_am_119, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_119), .B(
        b4_nUAi[992]), .C(b3_P_F_6_am_119), .Y(b6_2ZTGIf[330]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[330]), .B(
        b11_OFWNT9L_8tZ[46]), .C(b4_nUAi[991]), .D(b4_nUAi[990]), .Y(
        b3_P_F_6_am_119));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[330]), .B(
        b11_OFWNT9L_8tZ[46]), .C(b4_nUAi[990]), .D(b4_nUAi[991]), .Y(
        b3_P_F_6_bm_119));
    
endmodule


module b8_1LbcQDr1_x_107_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [269:269] mdiclink_reg;
input  [107:107] b11_OFWNT9L_8tZ;
input  [808:807] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[269]), .B(
        b11_OFWNT9L_8tZ[107]), .C(b4_nUAi[808]), .D(b4_nUAi[807]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[269]), .B(
        b11_OFWNT9L_8tZ[107]), .C(b4_nUAi[808]), .D(b4_nUAi[807]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_230_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [146:146] mdiclink_reg;
input  [230:230] b11_OFWNT9L_8tZ;
input  [440:438] b4_nUAi;
output [146:146] b6_2ZTGIf;

    wire b3_P_F_6_bm_36, b3_P_F_6_am_36, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_36), .B(
        b4_nUAi[440]), .C(b3_P_F_6_am_36), .Y(b6_2ZTGIf[146]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[146]), .B(
        b11_OFWNT9L_8tZ[230]), .C(b4_nUAi[439]), .D(b4_nUAi[438]), .Y(
        b3_P_F_6_am_36));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[146]), .B(
        b11_OFWNT9L_8tZ[230]), .C(b4_nUAi[438]), .D(b4_nUAi[439]), .Y(
        b3_P_F_6_bm_36));
    
endmodule


module b8_1LbcQDr1_x_198_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [178:178] mdiclink_reg;
input  [198:198] b11_OFWNT9L_8tZ;
input  [536:534] b4_nUAi;
output [178:178] b6_2ZTGIf;

    wire b3_P_F_6_bm_56, b3_P_F_6_am_56, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_56), .B(
        b4_nUAi[536]), .C(b3_P_F_6_am_56), .Y(b6_2ZTGIf[178]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[178]), .B(
        b11_OFWNT9L_8tZ[198]), .C(b4_nUAi[535]), .D(b4_nUAi[534]), .Y(
        b3_P_F_6_am_56));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[178]), .B(
        b11_OFWNT9L_8tZ[198]), .C(b4_nUAi[534]), .D(b4_nUAi[535]), .Y(
        b3_P_F_6_bm_56));
    
endmodule


module b8_1LbcQDr1_x_109_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [267:267] mdiclink_reg;
input  [109:109] b11_OFWNT9L_8tZ;
input  [802:801] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[267]), .B(
        b11_OFWNT9L_8tZ[109]), .C(b4_nUAi[802]), .D(b4_nUAi[801]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[267]), .B(
        b11_OFWNT9L_8tZ[109]), .C(b4_nUAi[802]), .D(b4_nUAi[801]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_223_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [153:153] mdiclink_reg;
input  [223:223] b11_OFWNT9L_8tZ;
input  [461:459] b4_nUAi;
output [153:153] b6_2ZTGIf;

    wire b3_P_F_6_bm_30, b3_P_F_6_am_30, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_30), .B(
        b4_nUAi[461]), .C(b3_P_F_6_am_30), .Y(b6_2ZTGIf[153]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[153]), .B(
        b11_OFWNT9L_8tZ[223]), .C(b4_nUAi[460]), .D(b4_nUAi[459]), .Y(
        b3_P_F_6_am_30));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[153]), .B(
        b11_OFWNT9L_8tZ[223]), .C(b4_nUAi[459]), .D(b4_nUAi[460]), .Y(
        b3_P_F_6_bm_30));
    
endmodule


module b8_1LbcQDr1_x_199_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [177:177] mdiclink_reg;
input  [199:199] b11_OFWNT9L_8tZ;
input  [533:531] b4_nUAi;
output [177:177] b6_2ZTGIf;

    wire b3_P_F_6_bm_57, b3_P_F_6_am_57, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_57), .B(
        b4_nUAi[533]), .C(b3_P_F_6_am_57), .Y(b6_2ZTGIf[177]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[177]), .B(
        b11_OFWNT9L_8tZ[199]), .C(b4_nUAi[532]), .D(b4_nUAi[531]), .Y(
        b3_P_F_6_am_57));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[177]), .B(
        b11_OFWNT9L_8tZ[199]), .C(b4_nUAi[531]), .D(b4_nUAi[532]), .Y(
        b3_P_F_6_bm_57));
    
endmodule


module b8_1LbcQDr1_x_352_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [24:24] mdiclink_reg;
input  [352:352] b11_OFWNT9L_8tZ;
input  [74:72] b4_nUAi;
output [24:24] b6_2ZTGIf;

    wire b3_P_F_6_bm_165, b3_P_F_6_am_165, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_165), .B(
        b4_nUAi[74]), .C(b3_P_F_6_am_165), .Y(b6_2ZTGIf[24]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[24]), .B(
        b11_OFWNT9L_8tZ[352]), .C(b4_nUAi[73]), .D(b4_nUAi[72]), .Y(
        b3_P_F_6_am_165));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[24]), .B(
        b11_OFWNT9L_8tZ[352]), .C(b4_nUAi[72]), .D(b4_nUAi[73]), .Y(
        b3_P_F_6_bm_165));
    
endmodule


module b8_1LbcQDr1_x_127_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [249:249] mdiclink_reg;
input  [127:127] b11_OFWNT9L_8tZ;
input  [749:747] b4_nUAi;
output [249:249] b6_2ZTGIf;

    wire b3_P_F_6_bm_224, b3_P_F_6_am_224, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_224), .B(
        b4_nUAi[749]), .C(b3_P_F_6_am_224), .Y(b6_2ZTGIf[249]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[249]), .B(
        b11_OFWNT9L_8tZ[127]), .C(b4_nUAi[748]), .D(b4_nUAi[747]), .Y(
        b3_P_F_6_am_224));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[249]), .B(
        b11_OFWNT9L_8tZ[127]), .C(b4_nUAi[747]), .D(b4_nUAi[748]), .Y(
        b3_P_F_6_bm_224));
    
endmodule


module b8_1LbcQDr1_x_158_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [218:218] mdiclink_reg;
input  [158:158] b11_OFWNT9L_8tZ;
input  [656:654] b4_nUAi;
output [218:218] b6_2ZTGIf;

    wire b3_P_F_6_bm_69, b3_P_F_6_am_69, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_69), .B(
        b4_nUAi[656]), .C(b3_P_F_6_am_69), .Y(b6_2ZTGIf[218]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[218]), .B(
        b11_OFWNT9L_8tZ[158]), .C(b4_nUAi[655]), .D(b4_nUAi[654]), .Y(
        b3_P_F_6_am_69));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[218]), .B(
        b11_OFWNT9L_8tZ[158]), .C(b4_nUAi[654]), .D(b4_nUAi[655]), .Y(
        b3_P_F_6_bm_69));
    
endmodule


module b8_1LbcQDr1_x_47_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [329:329] mdiclink_reg;
input  [47:47] b11_OFWNT9L_8tZ;
input  [989:987] b4_nUAi;
output [329:329] b6_2ZTGIf;

    wire b3_P_F_6_bm_120, b3_P_F_6_am_120, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_120), .B(
        b4_nUAi[989]), .C(b3_P_F_6_am_120), .Y(b6_2ZTGIf[329]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[329]), .B(
        b11_OFWNT9L_8tZ[47]), .C(b4_nUAi[988]), .D(b4_nUAi[987]), .Y(
        b3_P_F_6_am_120));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[329]), .B(
        b11_OFWNT9L_8tZ[47]), .C(b4_nUAi[987]), .D(b4_nUAi[988]), .Y(
        b3_P_F_6_bm_120));
    
endmodule


module b8_1LbcQDr1_x_354_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [22:22] mdiclink_reg;
input  [354:354] b11_OFWNT9L_8tZ;
input  [68:66] b4_nUAi;
output [22:22] b6_2ZTGIf;

    wire b3_P_F_6_bm_167, b3_P_F_6_am_167, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_167), .B(
        b4_nUAi[68]), .C(b3_P_F_6_am_167), .Y(b6_2ZTGIf[22]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[22]), .B(
        b11_OFWNT9L_8tZ[354]), .C(b4_nUAi[67]), .D(b4_nUAi[66]), .Y(
        b3_P_F_6_am_167));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[22]), .B(
        b11_OFWNT9L_8tZ[354]), .C(b4_nUAi[66]), .D(b4_nUAi[67]), .Y(
        b3_P_F_6_bm_167));
    
endmodule


module b8_1LbcQDr1_x_314_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [62:62] mdiclink_reg;
input  [314:314] b11_OFWNT9L_8tZ;
input  [187:186] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[62]), .B(
        b11_OFWNT9L_8tZ[314]), .C(b4_nUAi[187]), .D(b4_nUAi[186]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[62]), .B(
        b11_OFWNT9L_8tZ[314]), .C(b4_nUAi[187]), .D(b4_nUAi[186]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_168_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [208:208] mdiclink_reg;
input  [168:168] b11_OFWNT9L_8tZ;
input  [626:624] b4_nUAi;
output [208:208] b6_2ZTGIf;

    wire b3_P_F_6_bm_78, b3_P_F_6_am_78, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_78), .B(
        b4_nUAi[626]), .C(b3_P_F_6_am_78), .Y(b6_2ZTGIf[208]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[208]), .B(
        b11_OFWNT9L_8tZ[168]), .C(b4_nUAi[625]), .D(b4_nUAi[624]), .Y(
        b3_P_F_6_am_78));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[208]), .B(
        b11_OFWNT9L_8tZ[168]), .C(b4_nUAi[624]), .D(b4_nUAi[625]), .Y(
        b3_P_F_6_bm_78));
    
endmodule


module b8_1LbcQDr1_x_129_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [247:247] mdiclink_reg;
input  [129:129] b11_OFWNT9L_8tZ;
input  [743:741] b4_nUAi;
output [247:247] b6_2ZTGIf;

    wire b3_P_F_6_bm_226, b3_P_F_6_am_226, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_226), .B(
        b4_nUAi[743]), .C(b3_P_F_6_am_226), .Y(b6_2ZTGIf[247]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[247]), .B(
        b11_OFWNT9L_8tZ[129]), .C(b4_nUAi[742]), .D(b4_nUAi[741]), .Y(
        b3_P_F_6_am_226));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[247]), .B(
        b11_OFWNT9L_8tZ[129]), .C(b4_nUAi[741]), .D(b4_nUAi[742]), .Y(
        b3_P_F_6_bm_226));
    
endmodule


module b8_1LbcQDr1_x_206_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [170:170] mdiclink_reg;
input  [206:206] b11_OFWNT9L_8tZ;
input  [512:510] b4_nUAi;
output [170:170] b6_2ZTGIf;

    wire b3_P_F_6_bm_39, b3_P_F_6_am_39, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_39), .B(
        b4_nUAi[512]), .C(b3_P_F_6_am_39), .Y(b6_2ZTGIf[170]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[170]), .B(
        b11_OFWNT9L_8tZ[206]), .C(b4_nUAi[511]), .D(b4_nUAi[510]), .Y(
        b3_P_F_6_am_39));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[170]), .B(
        b11_OFWNT9L_8tZ[206]), .C(b4_nUAi[510]), .D(b4_nUAi[511]), .Y(
        b3_P_F_6_bm_39));
    
endmodule


module b8_1LbcQDr1_x_94_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [282:282] mdiclink_reg;
input  [94:94] b11_OFWNT9L_8tZ;
input  [848:846] b4_nUAi;
output [282:282] b6_2ZTGIf;

    wire b3_P_F_6_bm_89, b3_P_F_6_am_89, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_89), .B(
        b4_nUAi[848]), .C(b3_P_F_6_am_89), .Y(b6_2ZTGIf[282]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[282]), .B(
        b11_OFWNT9L_8tZ[94]), .C(b4_nUAi[847]), .D(b4_nUAi[846]), .Y(
        b3_P_F_6_am_89));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[282]), .B(
        b11_OFWNT9L_8tZ[94]), .C(b4_nUAi[846]), .D(b4_nUAi[847]), .Y(
        b3_P_F_6_bm_89));
    
endmodule


module b8_1LbcQDr1_x_1_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [375:375] mdiclink_reg;
input  [1:1] b11_OFWNT9L_8tZ;
input  [1127:1125] b4_nUAi;
output [375:375] b6_2ZTGIf;

    wire b3_P_F_6_bm_149, b3_P_F_6_am_149, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_149), .B(
        b4_nUAi[1127]), .C(b3_P_F_6_am_149), .Y(b6_2ZTGIf[375]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[375]), .B(
        b11_OFWNT9L_8tZ[1]), .C(b4_nUAi[1126]), .D(b4_nUAi[1125]), .Y(
        b3_P_F_6_am_149));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[375]), .B(
        b11_OFWNT9L_8tZ[1]), .C(b4_nUAi[1125]), .D(b4_nUAi[1126]), .Y(
        b3_P_F_6_bm_149));
    
endmodule


module b8_1LbcQDr1_x_335_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [41:41] mdiclink_reg;
input  [335:335] b11_OFWNT9L_8tZ;
input  [125:123] b4_nUAi;
output [41:41] b6_2ZTGIf;

    wire b3_P_F_6_bm_174, b3_P_F_6_am_174, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_174), .B(
        b4_nUAi[125]), .C(b3_P_F_6_am_174), .Y(b6_2ZTGIf[41]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[41]), .B(
        b11_OFWNT9L_8tZ[335]), .C(b4_nUAi[124]), .D(b4_nUAi[123]), .Y(
        b3_P_F_6_am_174));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[41]), .B(
        b11_OFWNT9L_8tZ[335]), .C(b4_nUAi[123]), .D(b4_nUAi[124]), .Y(
        b3_P_F_6_bm_174));
    
endmodule


module b8_1LbcQDr1_x_298_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [78:78] mdiclink_reg;
input  [298:298] b11_OFWNT9L_8tZ;
input  [235:234] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[78]), .B(
        b11_OFWNT9L_8tZ[298]), .C(b4_nUAi[235]), .D(b4_nUAi[234]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[78]), .B(
        b11_OFWNT9L_8tZ[298]), .C(b4_nUAi[235]), .D(b4_nUAi[234]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_358_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [18:18] mdiclink_reg;
input  [358:358] b11_OFWNT9L_8tZ;
input  [56:54] b4_nUAi;
output [18:18] b6_2ZTGIf;

    wire b3_P_F_6_bm_170, b3_P_F_6_am_170, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_170), .B(
        b4_nUAi[56]), .C(b3_P_F_6_am_170), .Y(b6_2ZTGIf[18]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[18]), .B(
        b11_OFWNT9L_8tZ[358]), .C(b4_nUAi[55]), .D(b4_nUAi[54]), .Y(
        b3_P_F_6_am_170));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[18]), .B(
        b11_OFWNT9L_8tZ[358]), .C(b4_nUAi[54]), .D(b4_nUAi[55]), .Y(
        b3_P_F_6_bm_170));
    
endmodule


module b8_1LbcQDr1_x_155_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [221:221] mdiclink_reg;
input  [155:155] b11_OFWNT9L_8tZ;
input  [664:663] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[221]), .B(
        b11_OFWNT9L_8tZ[155]), .C(b4_nUAi[664]), .D(b4_nUAi[663]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[221]), .B(
        b11_OFWNT9L_8tZ[155]), .C(b4_nUAi[664]), .D(b4_nUAi[663]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_62_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [314:314] mdiclink_reg;
input  [62:62] b11_OFWNT9L_8tZ;
input  [944:942] b4_nUAi;
output [314:314] b6_2ZTGIf;

    wire b3_P_F_6_bm_109, b3_P_F_6_am_109, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_109), .B(
        b4_nUAi[944]), .C(b3_P_F_6_am_109), .Y(b6_2ZTGIf[314]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[314]), .B(
        b11_OFWNT9L_8tZ[62]), .C(b4_nUAi[943]), .D(b4_nUAi[942]), .Y(
        b3_P_F_6_am_109));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[314]), .B(
        b11_OFWNT9L_8tZ[62]), .C(b4_nUAi[942]), .D(b4_nUAi[943]), .Y(
        b3_P_F_6_bm_109));
    
endmodule


module b8_1LbcQDr1_x_38_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [338:338] mdiclink_reg;
input  [38:38] b11_OFWNT9L_8tZ;
input  [1016:1014] b4_nUAi;
output [338:338] b6_2ZTGIf;

    wire b3_P_F_6_bm_136, b3_P_F_6_am_136, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_136), .B(
        b4_nUAi[1016]), .C(b3_P_F_6_am_136), .Y(b6_2ZTGIf[338]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[338]), .B(
        b11_OFWNT9L_8tZ[38]), .C(b4_nUAi[1015]), .D(b4_nUAi[1014]), .Y(
        b3_P_F_6_am_136));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[338]), .B(
        b11_OFWNT9L_8tZ[38]), .C(b4_nUAi[1014]), .D(b4_nUAi[1015]), .Y(
        b3_P_F_6_bm_136));
    
endmodule


module b8_1LbcQDr1_x_289_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [87:87] mdiclink_reg;
input  [289:289] b11_OFWNT9L_8tZ;
input  [263:261] b4_nUAi;
output [87:87] b6_2ZTGIf;

    wire b3_P_F_6_bm_206, b3_P_F_6_am_206, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_206), .B(
        b4_nUAi[263]), .C(b3_P_F_6_am_206), .Y(b6_2ZTGIf[87]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[87]), .B(
        b11_OFWNT9L_8tZ[289]), .C(b4_nUAi[262]), .D(b4_nUAi[261]), .Y(
        b3_P_F_6_am_206));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[87]), .B(
        b11_OFWNT9L_8tZ[289]), .C(b4_nUAi[261]), .D(b4_nUAi[262]), .Y(
        b3_P_F_6_bm_206));
    
endmodule


module b8_1LbcQDr1_x_336_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [40:40] mdiclink_reg;
input  [336:336] b11_OFWNT9L_8tZ;
input  [122:120] b4_nUAi;
output [40:40] b6_2ZTGIf;

    wire b3_P_F_6_bm_175, b3_P_F_6_am_175, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_175), .B(
        b4_nUAi[122]), .C(b3_P_F_6_am_175), .Y(b6_2ZTGIf[40]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[40]), .B(
        b11_OFWNT9L_8tZ[336]), .C(b4_nUAi[121]), .D(b4_nUAi[120]), .Y(
        b3_P_F_6_am_175));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[40]), .B(
        b11_OFWNT9L_8tZ[336]), .C(b4_nUAi[120]), .D(b4_nUAi[121]), .Y(
        b3_P_F_6_bm_175));
    
endmodule


module b8_1LbcQDr1_x_340_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [36:36] mdiclink_reg;
input  [340:340] b11_OFWNT9L_8tZ;
input  [110:108] b4_nUAi;
output [36:36] b6_2ZTGIf;

    wire b3_P_F_6_bm_178, b3_P_F_6_am_178, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_178), .B(
        b4_nUAi[110]), .C(b3_P_F_6_am_178), .Y(b6_2ZTGIf[36]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[36]), .B(
        b11_OFWNT9L_8tZ[340]), .C(b4_nUAi[109]), .D(b4_nUAi[108]), .Y(
        b3_P_F_6_am_178));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[36]), .B(
        b11_OFWNT9L_8tZ[340]), .C(b4_nUAi[108]), .D(b4_nUAi[109]), .Y(
        b3_P_F_6_bm_178));
    
endmodule


module b8_1LbcQDr1_x_166_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [210:210] mdiclink_reg;
input  [166:166] b11_OFWNT9L_8tZ;
input  [632:630] b4_nUAi;
output [210:210] b6_2ZTGIf;

    wire b3_P_F_6_bm_76, b3_P_F_6_am_76, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_76), .B(
        b4_nUAi[632]), .C(b3_P_F_6_am_76), .Y(b6_2ZTGIf[210]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[210]), .B(
        b11_OFWNT9L_8tZ[166]), .C(b4_nUAi[631]), .D(b4_nUAi[630]), .Y(
        b3_P_F_6_am_76));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[210]), .B(
        b11_OFWNT9L_8tZ[166]), .C(b4_nUAi[630]), .D(b4_nUAi[631]), .Y(
        b3_P_F_6_bm_76));
    
endmodule


module b8_1LbcQDr1_x_72_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [304:304] mdiclink_reg;
input  [72:72] b11_OFWNT9L_8tZ;
input  [914:912] b4_nUAi;
output [304:304] b6_2ZTGIf;

    wire b3_P_F_6_bm_118, b3_P_F_6_am_118, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_118), .B(
        b4_nUAi[914]), .C(b3_P_F_6_am_118), .Y(b6_2ZTGIf[304]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[304]), .B(
        b11_OFWNT9L_8tZ[72]), .C(b4_nUAi[913]), .D(b4_nUAi[912]), .Y(
        b3_P_F_6_am_118));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[304]), .B(
        b11_OFWNT9L_8tZ[72]), .C(b4_nUAi[912]), .D(b4_nUAi[913]), .Y(
        b3_P_F_6_bm_118));
    
endmodule


module b8_1LbcQDr1_x_318_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [58:58] mdiclink_reg;
input  [318:318] b11_OFWNT9L_8tZ;
input  [176:174] b4_nUAi;
output [58:58] b6_2ZTGIf;

    wire b3_P_F_6_bm_183, b3_P_F_6_am_183, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_183), .B(
        b4_nUAi[176]), .C(b3_P_F_6_am_183), .Y(b6_2ZTGIf[58]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[58]), .B(
        b11_OFWNT9L_8tZ[318]), .C(b4_nUAi[175]), .D(b4_nUAi[174]), .Y(
        b3_P_F_6_am_183));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[58]), .B(
        b11_OFWNT9L_8tZ[318]), .C(b4_nUAi[174]), .D(b4_nUAi[175]), .Y(
        b3_P_F_6_bm_183));
    
endmodule


module b8_1LbcQDr1_x_176_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [200:200] mdiclink_reg;
input  [176:176] b11_OFWNT9L_8tZ;
input  [602:600] b4_nUAi;
output [200:200] b6_2ZTGIf;

    wire b3_P_F_6_bm_61, b3_P_F_6_am_61, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_61), .B(
        b4_nUAi[602]), .C(b3_P_F_6_am_61), .Y(b6_2ZTGIf[200]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[200]), .B(
        b11_OFWNT9L_8tZ[176]), .C(b4_nUAi[601]), .D(b4_nUAi[600]), .Y(
        b3_P_F_6_am_61));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[200]), .B(
        b11_OFWNT9L_8tZ[176]), .C(b4_nUAi[600]), .D(b4_nUAi[601]), .Y(
        b3_P_F_6_bm_61));
    
endmodule


module b8_1LbcQDr1_x_205_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [171:171] mdiclink_reg;
input  [205:205] b11_OFWNT9L_8tZ;
input  [514:513] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[171]), .B(
        b11_OFWNT9L_8tZ[205]), .C(b4_nUAi[514]), .D(b4_nUAi[513]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[171]), .B(
        b11_OFWNT9L_8tZ[205]), .C(b4_nUAi[514]), .D(b4_nUAi[513]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_253_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [123:123] mdiclink_reg;
input  [253:253] b11_OFWNT9L_8tZ;
input  [370:369] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[123]), .B(
        b11_OFWNT9L_8tZ[253]), .C(b4_nUAi[370]), .D(b4_nUAi[369]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[123]), .B(
        b11_OFWNT9L_8tZ[253]), .C(b4_nUAi[370]), .D(b4_nUAi[369]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_66_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [310:310] mdiclink_reg;
input  [66:66] b11_OFWNT9L_8tZ;
input  [932:930] b4_nUAi;
output [310:310] b6_2ZTGIf;

    wire b3_P_F_6_bm_113, b3_P_F_6_am_113, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_113), .B(
        b4_nUAi[932]), .C(b3_P_F_6_am_113), .Y(b6_2ZTGIf[310]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[310]), .B(
        b11_OFWNT9L_8tZ[66]), .C(b4_nUAi[931]), .D(b4_nUAi[930]), .Y(
        b3_P_F_6_am_113));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[310]), .B(
        b11_OFWNT9L_8tZ[66]), .C(b4_nUAi[930]), .D(b4_nUAi[931]), .Y(
        b3_P_F_6_bm_113));
    
endmodule


module b8_1LbcQDr1_x_84_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [292:292] mdiclink_reg;
input  [84:84] b11_OFWNT9L_8tZ;
input  [878:876] b4_nUAi;
output [292:292] b6_2ZTGIf;

    wire b3_P_F_6_bm_104, b3_P_F_6_am_104, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_104), .B(
        b4_nUAi[878]), .C(b3_P_F_6_am_104), .Y(b6_2ZTGIf[292]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[292]), .B(
        b11_OFWNT9L_8tZ[84]), .C(b4_nUAi[877]), .D(b4_nUAi[876]), .Y(
        b3_P_F_6_am_104));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[292]), .B(
        b11_OFWNT9L_8tZ[84]), .C(b4_nUAi[876]), .D(b4_nUAi[877]), .Y(
        b3_P_F_6_bm_104));
    
endmodule


module b8_1LbcQDr1_x_76_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [300:300] mdiclink_reg;
input  [76:76] b11_OFWNT9L_8tZ;
input  [901:900] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[300]), .B(
        b11_OFWNT9L_8tZ[76]), .C(b4_nUAi[901]), .D(b4_nUAi[900]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[300]), .B(
        b11_OFWNT9L_8tZ[76]), .C(b4_nUAi[901]), .D(b4_nUAi[900]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_297_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [79:79] mdiclink_reg;
input  [297:297] b11_OFWNT9L_8tZ;
input  [238:237] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[79]), .B(
        b11_OFWNT9L_8tZ[297]), .C(b4_nUAi[238]), .D(b4_nUAi[237]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[79]), .B(
        b11_OFWNT9L_8tZ[297]), .C(b4_nUAi[238]), .D(b4_nUAi[237]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_357_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [19:19] mdiclink_reg;
input  [357:357] b11_OFWNT9L_8tZ;
input  [59:57] b4_nUAi;
output [19:19] b6_2ZTGIf;

    wire b3_P_F_6_bm_169, b3_P_F_6_am_169, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_169), .B(
        b4_nUAi[59]), .C(b3_P_F_6_am_169), .Y(b6_2ZTGIf[19]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[19]), .B(
        b11_OFWNT9L_8tZ[357]), .C(b4_nUAi[58]), .D(b4_nUAi[57]), .Y(
        b3_P_F_6_am_169));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[19]), .B(
        b11_OFWNT9L_8tZ[357]), .C(b4_nUAi[57]), .D(b4_nUAi[58]), .Y(
        b3_P_F_6_bm_169));
    
endmodule


module b8_1LbcQDr1_x_4_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [372:372] mdiclink_reg;
input  [4:4] b11_OFWNT9L_8tZ;
input  [1117:1116] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[372]), .B(
        b11_OFWNT9L_8tZ[4]), .C(b4_nUAi[1117]), .D(b4_nUAi[1116]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[372]), .B(
        b11_OFWNT9L_8tZ[4]), .C(b4_nUAi[1117]), .D(b4_nUAi[1116]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_110_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [266:266] mdiclink_reg;
input  [110:110] b11_OFWNT9L_8tZ;
input  [800:798] b4_nUAi;
output [266:266] b6_2ZTGIf;

    wire b3_P_F_6_bm_79, b3_P_F_6_am_79, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_79), .B(
        b4_nUAi[800]), .C(b3_P_F_6_am_79), .Y(b6_2ZTGIf[266]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[266]), .B(
        b11_OFWNT9L_8tZ[110]), .C(b4_nUAi[799]), .D(b4_nUAi[798]), .Y(
        b3_P_F_6_am_79));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[266]), .B(
        b11_OFWNT9L_8tZ[110]), .C(b4_nUAi[798]), .D(b4_nUAi[799]), .Y(
        b3_P_F_6_bm_79));
    
endmodule


module b8_1LbcQDr1_x_242_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [134:134] mdiclink_reg;
input  [242:242] b11_OFWNT9L_8tZ;
input  [404:402] b4_nUAi;
output [134:134] b6_2ZTGIf;

    wire b3_P_F_6_bm_23, b3_P_F_6_am_23, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_23), .B(
        b4_nUAi[404]), .C(b3_P_F_6_am_23), .Y(b6_2ZTGIf[134]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[134]), .B(
        b11_OFWNT9L_8tZ[242]), .C(b4_nUAi[403]), .D(b4_nUAi[402]), .Y(
        b3_P_F_6_am_23));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[134]), .B(
        b11_OFWNT9L_8tZ[242]), .C(b4_nUAi[402]), .D(b4_nUAi[403]), .Y(
        b3_P_F_6_bm_23));
    
endmodule


module b8_1LbcQDr1_x_317_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [59:59] mdiclink_reg;
input  [317:317] b11_OFWNT9L_8tZ;
input  [178:177] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[59]), .B(
        b11_OFWNT9L_8tZ[317]), .C(b4_nUAi[178]), .D(b4_nUAi[177]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[59]), .B(
        b11_OFWNT9L_8tZ[317]), .C(b4_nUAi[178]), .D(b4_nUAi[177]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_372_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [4:4] mdiclink_reg;
input  [372:372] b11_OFWNT9L_8tZ;
input  [14:12] b4_nUAi;
output [4:4] b6_2ZTGIf;

    wire b3_P_F_6_bm_158, b3_P_F_6_am_158, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_158), .B(
        b4_nUAi[14]), .C(b3_P_F_6_am_158), .Y(b6_2ZTGIf[4]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[4]), .B(
        b11_OFWNT9L_8tZ[372]), .C(b4_nUAi[13]), .D(b4_nUAi[12]), .Y(
        b3_P_F_6_am_158));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[4]), .B(
        b11_OFWNT9L_8tZ[372]), .C(b4_nUAi[12]), .D(b4_nUAi[13]), .Y(
        b3_P_F_6_bm_158));
    
endmodule


module b8_1LbcQDr1_x_240_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [136:136] mdiclink_reg;
input  [240:240] b11_OFWNT9L_8tZ;
input  [410:408] b4_nUAi;
output [136:136] b6_2ZTGIf;

    wire b3_P_F_6_bm_21, b3_P_F_6_am_21, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_21), .B(
        b4_nUAi[410]), .C(b3_P_F_6_am_21), .Y(b6_2ZTGIf[136]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[136]), .B(
        b11_OFWNT9L_8tZ[240]), .C(b4_nUAi[409]), .D(b4_nUAi[408]), .Y(
        b3_P_F_6_am_21));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[136]), .B(
        b11_OFWNT9L_8tZ[240]), .C(b4_nUAi[408]), .D(b4_nUAi[409]), .Y(
        b3_P_F_6_bm_21));
    
endmodule


module b8_1LbcQDr1_x_122_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [254:254] mdiclink_reg;
input  [122:122] b11_OFWNT9L_8tZ;
input  [763:762] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[254]), .B(
        b11_OFWNT9L_8tZ[122]), .C(b4_nUAi[763]), .D(b4_nUAi[762]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[254]), .B(
        b11_OFWNT9L_8tZ[122]), .C(b4_nUAi[763]), .D(b4_nUAi[762]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_130_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [246:246] mdiclink_reg;
input  [130:130] b11_OFWNT9L_8tZ;
input  [740:738] b4_nUAi;
output [246:246] b6_2ZTGIf;

    wire b3_P_F_6_bm_227, b3_P_F_6_am_227, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_227), .B(
        b4_nUAi[740]), .C(b3_P_F_6_am_227), .Y(b6_2ZTGIf[246]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[246]), .B(
        b11_OFWNT9L_8tZ[130]), .C(b4_nUAi[739]), .D(b4_nUAi[738]), .Y(
        b3_P_F_6_am_227));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[246]), .B(
        b11_OFWNT9L_8tZ[130]), .C(b4_nUAi[738]), .D(b4_nUAi[739]), .Y(
        b3_P_F_6_bm_227));
    
endmodule


module b8_1LbcQDr1_x_137_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [239:239] mdiclink_reg;
input  [137:137] b11_OFWNT9L_8tZ;
input  [718:717] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[239]), .B(
        b11_OFWNT9L_8tZ[137]), .C(b4_nUAi[718]), .D(b4_nUAi[717]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[239]), .B(
        b11_OFWNT9L_8tZ[137]), .C(b4_nUAi[718]), .D(b4_nUAi[717]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_93_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [283:283] mdiclink_reg;
input  [93:93] b11_OFWNT9L_8tZ;
input  [850:849] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[283]), .B(
        b11_OFWNT9L_8tZ[93]), .C(b4_nUAi[850]), .D(b4_nUAi[849]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[283]), .B(
        b11_OFWNT9L_8tZ[93]), .C(b4_nUAi[850]), .D(b4_nUAi[849]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_20_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [356:356] mdiclink_reg;
input  [20:20] b11_OFWNT9L_8tZ;
input  [1070:1068] b4_nUAi;
output [356:356] b6_2ZTGIf;

    wire b3_P_F_6_bm_144, b3_P_F_6_am_144, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_144), .B(
        b4_nUAi[1070]), .C(b3_P_F_6_am_144), .Y(b6_2ZTGIf[356]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[356]), .B(
        b11_OFWNT9L_8tZ[20]), .C(b4_nUAi[1069]), .D(b4_nUAi[1068]), .Y(
        b3_P_F_6_am_144));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[356]), .B(
        b11_OFWNT9L_8tZ[20]), .C(b4_nUAi[1068]), .D(b4_nUAi[1069]), .Y(
        b3_P_F_6_bm_144));
    
endmodule


module b8_1LbcQDr1_x_139_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [237:237] mdiclink_reg;
input  [139:139] b11_OFWNT9L_8tZ;
input  [712:711] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[237]), .B(
        b11_OFWNT9L_8tZ[139]), .C(b4_nUAi[712]), .D(b4_nUAi[711]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[237]), .B(
        b11_OFWNT9L_8tZ[139]), .C(b4_nUAi[712]), .D(b4_nUAi[711]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_58_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [318:318] mdiclink_reg;
input  [58:58] b11_OFWNT9L_8tZ;
input  [955:954] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[318]), .B(
        b11_OFWNT9L_8tZ[58]), .C(b4_nUAi[955]), .D(b4_nUAi[954]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[318]), .B(
        b11_OFWNT9L_8tZ[58]), .C(b4_nUAi[955]), .D(b4_nUAi[954]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_68_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [308:308] mdiclink_reg;
input  [68:68] b11_OFWNT9L_8tZ;
input  [926:924] b4_nUAi;
output [308:308] b6_2ZTGIf;

    wire b3_P_F_6_bm_114, b3_P_F_6_am_114, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_114), .B(
        b4_nUAi[926]), .C(b3_P_F_6_am_114), .Y(b6_2ZTGIf[308]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[308]), .B(
        b11_OFWNT9L_8tZ[68]), .C(b4_nUAi[925]), .D(b4_nUAi[924]), .Y(
        b3_P_F_6_am_114));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[308]), .B(
        b11_OFWNT9L_8tZ[68]), .C(b4_nUAi[924]), .D(b4_nUAi[925]), .Y(
        b3_P_F_6_bm_114));
    
endmodule


module b8_1LbcQDr1_x_349_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [27:27] mdiclink_reg;
input  [349:349] b11_OFWNT9L_8tZ;
input  [82:81] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[27]), .B(
        b11_OFWNT9L_8tZ[349]), .C(b4_nUAi[82]), .D(b4_nUAi[81]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[27]), .B(
        b11_OFWNT9L_8tZ[349]), .C(b4_nUAi[82]), .D(b4_nUAi[81]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_83_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [293:293] mdiclink_reg;
input  [83:83] b11_OFWNT9L_8tZ;
input  [880:879] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[293]), .B(
        b11_OFWNT9L_8tZ[83]), .C(b4_nUAi[880]), .D(b4_nUAi[879]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[293]), .B(
        b11_OFWNT9L_8tZ[83]), .C(b4_nUAi[880]), .D(b4_nUAi[879]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_309_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [67:67] mdiclink_reg;
input  [309:309] b11_OFWNT9L_8tZ;
input  [203:201] b4_nUAi;
output [67:67] b6_2ZTGIf;

    wire b3_P_F_6_bm_199, b3_P_F_6_am_199, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_199), .B(
        b4_nUAi[203]), .C(b3_P_F_6_am_199), .Y(b6_2ZTGIf[67]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[67]), .B(
        b11_OFWNT9L_8tZ[309]), .C(b4_nUAi[202]), .D(b4_nUAi[201]), .Y(
        b3_P_F_6_am_199));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[67]), .B(
        b11_OFWNT9L_8tZ[309]), .C(b4_nUAi[201]), .D(b4_nUAi[202]), .Y(
        b3_P_F_6_bm_199));
    
endmodule


module b8_1LbcQDr1_x_152_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [224:224] mdiclink_reg;
input  [152:152] b11_OFWNT9L_8tZ;
input  [674:672] b4_nUAi;
output [224:224] b6_2ZTGIf;

    wire b3_P_F_6_bm_222, b3_P_F_6_am_222, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_222), .B(
        b4_nUAi[674]), .C(b3_P_F_6_am_222), .Y(b6_2ZTGIf[224]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[224]), .B(
        b11_OFWNT9L_8tZ[152]), .C(b4_nUAi[673]), .D(b4_nUAi[672]), .Y(
        b3_P_F_6_am_222));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[224]), .B(
        b11_OFWNT9L_8tZ[152]), .C(b4_nUAi[672]), .D(b4_nUAi[673]), .Y(
        b3_P_F_6_bm_222));
    
endmodule


module b8_1LbcQDr1_x_19_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [357:357] mdiclink_reg;
input  [19:19] b11_OFWNT9L_8tZ;
input  [1072:1071] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[357]), .B(
        b11_OFWNT9L_8tZ[19]), .C(b4_nUAi[1072]), .D(b4_nUAi[1071]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[357]), .B(
        b11_OFWNT9L_8tZ[19]), .C(b4_nUAi[1072]), .D(b4_nUAi[1071]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_262_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [114:114] mdiclink_reg;
input  [262:262] b11_OFWNT9L_8tZ;
input  [344:342] b4_nUAi;
output [114:114] b6_2ZTGIf;

    wire b3_P_F_6_bm_16, b3_P_F_6_am_16, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_16), .B(
        b4_nUAi[344]), .C(b3_P_F_6_am_16), .Y(b6_2ZTGIf[114]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[114]), .B(
        b11_OFWNT9L_8tZ[262]), .C(b4_nUAi[343]), .D(b4_nUAi[342]), .Y(
        b3_P_F_6_am_16));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[114]), .B(
        b11_OFWNT9L_8tZ[262]), .C(b4_nUAi[342]), .D(b4_nUAi[343]), .Y(
        b3_P_F_6_bm_16));
    
endmodule


module b8_1LbcQDr1_x_88_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [288:288] mdiclink_reg;
input  [88:88] b11_OFWNT9L_8tZ;
input  [866:864] b4_nUAi;
output [288:288] b6_2ZTGIf;

    wire b3_P_F_6_bm_108, b3_P_F_6_am_108, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_108), .B(
        b4_nUAi[866]), .C(b3_P_F_6_am_108), .Y(b6_2ZTGIf[288]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[288]), .B(
        b11_OFWNT9L_8tZ[88]), .C(b4_nUAi[865]), .D(b4_nUAi[864]), .Y(
        b3_P_F_6_am_108));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[288]), .B(
        b11_OFWNT9L_8tZ[88]), .C(b4_nUAi[864]), .D(b4_nUAi[865]), .Y(
        b3_P_F_6_bm_108));
    
endmodule


module b8_1LbcQDr1_x_280_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [96:96] mdiclink_reg;
input  [280:280] b11_OFWNT9L_8tZ;
input  [290:288] b4_nUAi;
output [96:96] b6_2ZTGIf;

    wire b3_P_F_6_bm_8, b3_P_F_6_am_8, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_8), .B(
        b4_nUAi[290]), .C(b3_P_F_6_am_8), .Y(b6_2ZTGIf[96]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[96]), .B(
        b11_OFWNT9L_8tZ[280]), .C(b4_nUAi[289]), .D(b4_nUAi[288]), .Y(
        b3_P_F_6_am_8));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[96]), .B(
        b11_OFWNT9L_8tZ[280]), .C(b4_nUAi[288]), .D(b4_nUAi[289]), .Y(
        b3_P_F_6_bm_8));
    
endmodule


module b8_1LbcQDr1_x_260_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [116:116] mdiclink_reg;
input  [260:260] b11_OFWNT9L_8tZ;
input  [350:348] b4_nUAi;
output [116:116] b6_2ZTGIf;

    wire b3_P_F_6_bm_14, b3_P_F_6_am_14, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_14), .B(
        b4_nUAi[350]), .C(b3_P_F_6_am_14), .Y(b6_2ZTGIf[116]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[116]), .B(
        b11_OFWNT9L_8tZ[260]), .C(b4_nUAi[349]), .D(b4_nUAi[348]), .Y(
        b3_P_F_6_am_14));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[116]), .B(
        b11_OFWNT9L_8tZ[260]), .C(b4_nUAi[348]), .D(b4_nUAi[349]), .Y(
        b3_P_F_6_bm_14));
    
endmodule


module b8_1LbcQDr1_x_105_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [271:271] mdiclink_reg;
input  [105:105] b11_OFWNT9L_8tZ;
input  [814:813] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[271]), .B(
        b11_OFWNT9L_8tZ[105]), .C(b4_nUAi[814]), .D(b4_nUAi[813]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[271]), .B(
        b11_OFWNT9L_8tZ[105]), .C(b4_nUAi[814]), .D(b4_nUAi[813]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_272_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [104:104] mdiclink_reg;
input  [272:272] b11_OFWNT9L_8tZ;
input  [314:312] b4_nUAi;
output [104:104] b6_2ZTGIf;

    wire b3_P_F_6_bm_1, b3_P_F_6_am_1, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_1), .B(
        b4_nUAi[314]), .C(b3_P_F_6_am_1), .Y(b6_2ZTGIf[104]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[104]), .B(
        b11_OFWNT9L_8tZ[272]), .C(b4_nUAi[313]), .D(b4_nUAi[312]), .Y(
        b3_P_F_6_am_1));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[104]), .B(
        b11_OFWNT9L_8tZ[272]), .C(b4_nUAi[312]), .D(b4_nUAi[313]), .Y(
        b3_P_F_6_bm_1));
    
endmodule


module b8_1LbcQDr1_x_343_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [33:33] mdiclink_reg;
input  [343:343] b11_OFWNT9L_8tZ;
input  [101:99] b4_nUAi;
output [33:33] b6_2ZTGIf;

    wire b3_P_F_6_bm_181, b3_P_F_6_am_181, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_181), .B(
        b4_nUAi[101]), .C(b3_P_F_6_am_181), .Y(b6_2ZTGIf[33]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[33]), .B(
        b11_OFWNT9L_8tZ[343]), .C(b4_nUAi[100]), .D(b4_nUAi[99]), .Y(
        b3_P_F_6_am_181));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[33]), .B(
        b11_OFWNT9L_8tZ[343]), .C(b4_nUAi[99]), .D(b4_nUAi[100]), .Y(
        b3_P_F_6_bm_181));
    
endmodule


module b8_1LbcQDr1_x_270_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [106:106] mdiclink_reg;
input  [270:270] b11_OFWNT9L_8tZ;
input  [320:318] b4_nUAi;
output [106:106] b6_2ZTGIf;

    wire b3_P_F_6_bm_net_1, b3_P_F_6_am_net_1, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_net_1), .B(
        b4_nUAi[320]), .C(b3_P_F_6_am_net_1), .Y(b6_2ZTGIf[106]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[106]), .B(
        b11_OFWNT9L_8tZ[270]), .C(b4_nUAi[319]), .D(b4_nUAi[318]), .Y(
        b3_P_F_6_am_net_1));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[106]), .B(
        b11_OFWNT9L_8tZ[270]), .C(b4_nUAi[318]), .D(b4_nUAi[319]), .Y(
        b3_P_F_6_bm_net_1));
    
endmodule


module b8_1LbcQDr1_x_50_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [326:326] mdiclink_reg;
input  [50:50] b11_OFWNT9L_8tZ;
input  [980:978] b4_nUAi;
output [326:326] b6_2ZTGIf;

    wire b3_P_F_6_bm_123, b3_P_F_6_am_123, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_123), .B(
        b4_nUAi[980]), .C(b3_P_F_6_am_123), .Y(b6_2ZTGIf[326]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[326]), .B(
        b11_OFWNT9L_8tZ[50]), .C(b4_nUAi[979]), .D(b4_nUAi[978]), .Y(
        b3_P_F_6_am_123));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[326]), .B(
        b11_OFWNT9L_8tZ[50]), .C(b4_nUAi[978]), .D(b4_nUAi[979]), .Y(
        b3_P_F_6_bm_123));
    
endmodule


module b8_1LbcQDr1_x_124_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [252:252] mdiclink_reg;
input  [124:124] b11_OFWNT9L_8tZ;
input  [757:756] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[252]), .B(
        b11_OFWNT9L_8tZ[124]), .C(b4_nUAi[757]), .D(b4_nUAi[756]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[252]), .B(
        b11_OFWNT9L_8tZ[124]), .C(b4_nUAi[757]), .D(b4_nUAi[756]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_157_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [219:219] mdiclink_reg;
input  [157:157] b11_OFWNT9L_8tZ;
input  [658:657] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[219]), .B(
        b11_OFWNT9L_8tZ[157]), .C(b4_nUAi[658]), .D(b4_nUAi[657]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[219]), .B(
        b11_OFWNT9L_8tZ[157]), .C(b4_nUAi[658]), .D(b4_nUAi[657]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_203_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [173:173] mdiclink_reg;
input  [203:203] b11_OFWNT9L_8tZ;
input  [520:519] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[173]), .B(
        b11_OFWNT9L_8tZ[203]), .C(b4_nUAi[520]), .D(b4_nUAi[519]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[173]), .B(
        b11_OFWNT9L_8tZ[203]), .C(b4_nUAi[520]), .D(b4_nUAi[519]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_328_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [48:48] mdiclink_reg;
input  [328:328] b11_OFWNT9L_8tZ;
input  [146:144] b4_nUAi;
output [48:48] b6_2ZTGIf;

    wire b3_P_F_6_bm_192, b3_P_F_6_am_192, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_192), .B(
        b4_nUAi[146]), .C(b3_P_F_6_am_192), .Y(b6_2ZTGIf[48]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[48]), .B(
        b11_OFWNT9L_8tZ[328]), .C(b4_nUAi[145]), .D(b4_nUAi[144]), .Y(
        b3_P_F_6_am_192));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[48]), .B(
        b11_OFWNT9L_8tZ[328]), .C(b4_nUAi[144]), .D(b4_nUAi[145]), .Y(
        b3_P_F_6_bm_192));
    
endmodule


module b8_1LbcQDr1_x_301_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [75:75] mdiclink_reg;
input  [301:301] b11_OFWNT9L_8tZ;
input  [226:225] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[75]), .B(
        b11_OFWNT9L_8tZ[301]), .C(b4_nUAi[226]), .D(b4_nUAi[225]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[75]), .B(
        b11_OFWNT9L_8tZ[301]), .C(b4_nUAi[226]), .D(b4_nUAi[225]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_361_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [15:15] mdiclink_reg;
input  [361:361] b11_OFWNT9L_8tZ;
input  [46:45] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[15]), .B(
        b11_OFWNT9L_8tZ[361]), .C(b4_nUAi[46]), .D(b4_nUAi[45]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[15]), .B(
        b11_OFWNT9L_8tZ[361]), .C(b4_nUAi[46]), .D(b4_nUAi[45]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_78_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [298:298] mdiclink_reg;
input  [78:78] b11_OFWNT9L_8tZ;
input  [896:894] b4_nUAi;
output [298:298] b6_2ZTGIf;

    wire b3_P_F_6_bm_99, b3_P_F_6_am_99, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_99), .B(
        b4_nUAi[896]), .C(b3_P_F_6_am_99), .Y(b6_2ZTGIf[298]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[298]), .B(
        b11_OFWNT9L_8tZ[78]), .C(b4_nUAi[895]), .D(b4_nUAi[894]), .Y(
        b3_P_F_6_am_99));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[298]), .B(
        b11_OFWNT9L_8tZ[78]), .C(b4_nUAi[894]), .D(b4_nUAi[895]), .Y(
        b3_P_F_6_bm_99));
    
endmodule


module b8_1LbcQDr1_x_167_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [209:209] mdiclink_reg;
input  [167:167] b11_OFWNT9L_8tZ;
input  [629:627] b4_nUAi;
output [209:209] b6_2ZTGIf;

    wire b3_P_F_6_bm_77, b3_P_F_6_am_77, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_77), .B(
        b4_nUAi[629]), .C(b3_P_F_6_am_77), .Y(b6_2ZTGIf[209]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[209]), .B(
        b11_OFWNT9L_8tZ[167]), .C(b4_nUAi[628]), .D(b4_nUAi[627]), .Y(
        b3_P_F_6_am_77));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[209]), .B(
        b11_OFWNT9L_8tZ[167]), .C(b4_nUAi[627]), .D(b4_nUAi[628]), .Y(
        b3_P_F_6_bm_77));
    
endmodule


module b8_1LbcQDr1_x_159_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [217:217] mdiclink_reg;
input  [159:159] b11_OFWNT9L_8tZ;
input  [653:651] b4_nUAi;
output [217:217] b6_2ZTGIf;

    wire b3_P_F_6_bm_70, b3_P_F_6_am_70, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_70), .B(
        b4_nUAi[653]), .C(b3_P_F_6_am_70), .Y(b6_2ZTGIf[217]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[217]), .B(
        b11_OFWNT9L_8tZ[159]), .C(b4_nUAi[652]), .D(b4_nUAi[651]), .Y(
        b3_P_F_6_am_70));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[217]), .B(
        b11_OFWNT9L_8tZ[159]), .C(b4_nUAi[651]), .D(b4_nUAi[652]), .Y(
        b3_P_F_6_bm_70));
    
endmodule


module b8_1LbcQDr1_x_369_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [7:7] mdiclink_reg;
input  [369:369] b11_OFWNT9L_8tZ;
input  [23:21] b4_nUAi;
output [7:7] b6_2ZTGIf;

    wire b3_P_F_6_bm_156, b3_P_F_6_am_156, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_156), .B(
        b4_nUAi[23]), .C(b3_P_F_6_am_156), .Y(b6_2ZTGIf[7]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[7]), .B(
        b11_OFWNT9L_8tZ[369]), .C(b4_nUAi[22]), .D(b4_nUAi[21]), .Y(
        b3_P_F_6_am_156));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[7]), .B(
        b11_OFWNT9L_8tZ[369]), .C(b4_nUAi[21]), .D(b4_nUAi[22]), .Y(
        b3_P_F_6_bm_156));
    
endmodule


module b8_1LbcQDr1_x_96_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [280:280] mdiclink_reg;
input  [96:96] b11_OFWNT9L_8tZ;
input  [842:840] b4_nUAi;
output [280:280] b6_2ZTGIf;

    wire b3_P_F_6_bm_91, b3_P_F_6_am_91, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_91), .B(
        b4_nUAi[842]), .C(b3_P_F_6_am_91), .Y(b6_2ZTGIf[280]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[280]), .B(
        b11_OFWNT9L_8tZ[96]), .C(b4_nUAi[841]), .D(b4_nUAi[840]), .Y(
        b3_P_F_6_am_91));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[280]), .B(
        b11_OFWNT9L_8tZ[96]), .C(b4_nUAi[840]), .D(b4_nUAi[841]), .Y(
        b3_P_F_6_bm_91));
    
endmodule


module b8_1LbcQDr1_x_140_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [236:236] mdiclink_reg;
input  [140:140] b11_OFWNT9L_8tZ;
input  [709:708] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[236]), .B(
        b11_OFWNT9L_8tZ[140]), .C(b4_nUAi[709]), .D(b4_nUAi[708]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[236]), .B(
        b11_OFWNT9L_8tZ[140]), .C(b4_nUAi[709]), .D(b4_nUAi[708]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_13_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [363:363] mdiclink_reg;
input  [13:13] b11_OFWNT9L_8tZ;
input  [1090:1089] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[363]), .B(
        b11_OFWNT9L_8tZ[13]), .C(b4_nUAi[1090]), .D(b4_nUAi[1089]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[363]), .B(
        b11_OFWNT9L_8tZ[13]), .C(b4_nUAi[1090]), .D(b4_nUAi[1089]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_169_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [207:207] mdiclink_reg;
input  [169:169] b11_OFWNT9L_8tZ;
input  [622:621] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[207]), .B(
        b11_OFWNT9L_8tZ[169]), .C(b4_nUAi[622]), .D(b4_nUAi[621]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[207]), .B(
        b11_OFWNT9L_8tZ[169]), .C(b4_nUAi[622]), .D(b4_nUAi[621]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_321_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [55:55] mdiclink_reg;
input  [321:321] b11_OFWNT9L_8tZ;
input  [167:165] b4_nUAi;
output [55:55] b6_2ZTGIf;

    wire b3_P_F_6_bm_186, b3_P_F_6_am_186, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_186), .B(
        b4_nUAi[167]), .C(b3_P_F_6_am_186), .Y(b6_2ZTGIf[55]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[55]), .B(
        b11_OFWNT9L_8tZ[321]), .C(b4_nUAi[166]), .D(b4_nUAi[165]), .Y(
        b3_P_F_6_am_186));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[55]), .B(
        b11_OFWNT9L_8tZ[321]), .C(b4_nUAi[165]), .D(b4_nUAi[166]), .Y(
        b3_P_F_6_bm_186));
    
endmodule


module b8_1LbcQDr1_x_49_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [327:327] mdiclink_reg;
input  [49:49] b11_OFWNT9L_8tZ;
input  [983:981] b4_nUAi;
output [327:327] b6_2ZTGIf;

    wire b3_P_F_6_bm_122, b3_P_F_6_am_122, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_122), .B(
        b4_nUAi[983]), .C(b3_P_F_6_am_122), .Y(b6_2ZTGIf[327]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[327]), .B(
        b11_OFWNT9L_8tZ[49]), .C(b4_nUAi[982]), .D(b4_nUAi[981]), .Y(
        b3_P_F_6_am_122));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[327]), .B(
        b11_OFWNT9L_8tZ[49]), .C(b4_nUAi[981]), .D(b4_nUAi[982]), .Y(
        b3_P_F_6_bm_122));
    
endmodule


module b8_1LbcQDr1_x_327_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [49:49] mdiclink_reg;
input  [327:327] b11_OFWNT9L_8tZ;
input  [149:147] b4_nUAi;
output [49:49] b6_2ZTGIf;

    wire b3_P_F_6_bm_191, b3_P_F_6_am_191, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_191), .B(
        b4_nUAi[149]), .C(b3_P_F_6_am_191), .Y(b6_2ZTGIf[49]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[49]), .B(
        b11_OFWNT9L_8tZ[327]), .C(b4_nUAi[148]), .D(b4_nUAi[147]), .Y(
        b3_P_F_6_am_191));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[49]), .B(
        b11_OFWNT9L_8tZ[327]), .C(b4_nUAi[147]), .D(b4_nUAi[148]), .Y(
        b3_P_F_6_bm_191));
    
endmodule


module b8_1LbcQDr1_x_33_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [343:343] mdiclink_reg;
input  [33:33] b11_OFWNT9L_8tZ;
input  [1031:1029] b4_nUAi;
output [343:343] b6_2ZTGIf;

    wire b3_P_F_6_bm_132, b3_P_F_6_am_132, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_132), .B(
        b4_nUAi[1031]), .C(b3_P_F_6_am_132), .Y(b6_2ZTGIf[343]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[343]), .B(
        b11_OFWNT9L_8tZ[33]), .C(b4_nUAi[1030]), .D(b4_nUAi[1029]), .Y(
        b3_P_F_6_am_132));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[343]), .B(
        b11_OFWNT9L_8tZ[33]), .C(b4_nUAi[1029]), .D(b4_nUAi[1030]), .Y(
        b3_P_F_6_bm_132));
    
endmodule


module b8_1LbcQDr1_x_25_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [351:351] mdiclink_reg;
input  [25:25] b11_OFWNT9L_8tZ;
input  [1054:1053] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[351]), .B(
        b11_OFWNT9L_8tZ[25]), .C(b4_nUAi[1054]), .D(b4_nUAi[1053]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[351]), .B(
        b11_OFWNT9L_8tZ[25]), .C(b4_nUAi[1054]), .D(b4_nUAi[1053]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_86_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [290:290] mdiclink_reg;
input  [86:86] b11_OFWNT9L_8tZ;
input  [872:870] b4_nUAi;
output [290:290] b6_2ZTGIf;

    wire b3_P_F_6_bm_106, b3_P_F_6_am_106, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_106), .B(
        b4_nUAi[872]), .C(b3_P_F_6_am_106), .Y(b6_2ZTGIf[290]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[290]), .B(
        b11_OFWNT9L_8tZ[86]), .C(b4_nUAi[871]), .D(b4_nUAi[870]), .Y(
        b3_P_F_6_am_106));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[290]), .B(
        b11_OFWNT9L_8tZ[86]), .C(b4_nUAi[870]), .D(b4_nUAi[871]), .Y(
        b3_P_F_6_bm_106));
    
endmodule


module b8_1LbcQDr1_x_332_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [44:44] mdiclink_reg;
input  [332:332] b11_OFWNT9L_8tZ;
input  [133:132] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[44]), .B(
        b11_OFWNT9L_8tZ[332]), .C(b4_nUAi[133]), .D(b4_nUAi[132]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[44]), .B(
        b11_OFWNT9L_8tZ[332]), .C(b4_nUAi[133]), .D(b4_nUAi[132]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_154_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [222:222] mdiclink_reg;
input  [154:154] b11_OFWNT9L_8tZ;
input  [667:666] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[222]), .B(
        b11_OFWNT9L_8tZ[154]), .C(b4_nUAi[667]), .D(b4_nUAi[666]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[222]), .B(
        b11_OFWNT9L_8tZ[154]), .C(b4_nUAi[667]), .D(b4_nUAi[666]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_345_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [31:31] mdiclink_reg;
input  [345:345] b11_OFWNT9L_8tZ;
input  [94:93] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[31]), .B(
        b11_OFWNT9L_8tZ[345]), .C(b4_nUAi[94]), .D(b4_nUAi[93]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[31]), .B(
        b11_OFWNT9L_8tZ[345]), .C(b4_nUAi[94]), .D(b4_nUAi[93]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_111_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [265:265] mdiclink_reg;
input  [111:111] b11_OFWNT9L_8tZ;
input  [797:795] b4_nUAi;
output [265:265] b6_2ZTGIf;

    wire b3_P_F_6_bm_80, b3_P_F_6_am_80, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_80), .B(
        b4_nUAi[797]), .C(b3_P_F_6_am_80), .Y(b6_2ZTGIf[265]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[265]), .B(
        b11_OFWNT9L_8tZ[111]), .C(b4_nUAi[796]), .D(b4_nUAi[795]), .Y(
        b3_P_F_6_am_80));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[265]), .B(
        b11_OFWNT9L_8tZ[111]), .C(b4_nUAi[795]), .D(b4_nUAi[796]), .Y(
        b3_P_F_6_bm_80));
    
endmodule


module b8_1LbcQDr1_x_304_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [72:72] mdiclink_reg;
input  [304:304] b11_OFWNT9L_8tZ;
input  [218:216] b4_nUAi;
output [72:72] b6_2ZTGIf;

    wire b3_P_F_6_bm_195, b3_P_F_6_am_195, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_195), .B(
        b4_nUAi[218]), .C(b3_P_F_6_am_195), .Y(b6_2ZTGIf[72]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[72]), .B(
        b11_OFWNT9L_8tZ[304]), .C(b4_nUAi[217]), .D(b4_nUAi[216]), .Y(
        b3_P_F_6_am_195));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[72]), .B(
        b11_OFWNT9L_8tZ[304]), .C(b4_nUAi[216]), .D(b4_nUAi[217]), .Y(
        b3_P_F_6_bm_195));
    
endmodule


module b8_1LbcQDr1_x_364_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [12:12] mdiclink_reg;
input  [364:364] b11_OFWNT9L_8tZ;
input  [37:36] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[12]), .B(
        b11_OFWNT9L_8tZ[364]), .C(b4_nUAi[37]), .D(b4_nUAi[36]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[12]), .B(
        b11_OFWNT9L_8tZ[364]), .C(b4_nUAi[37]), .D(b4_nUAi[36]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_346_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [30:30] mdiclink_reg;
input  [346:346] b11_OFWNT9L_8tZ;
input  [91:90] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[30]), .B(
        b11_OFWNT9L_8tZ[346]), .C(b4_nUAi[91]), .D(b4_nUAi[90]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[30]), .B(
        b11_OFWNT9L_8tZ[346]), .C(b4_nUAi[91]), .D(b4_nUAi[90]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_214_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [162:162] mdiclink_reg;
input  [214:214] b11_OFWNT9L_8tZ;
input  [488:486] b4_nUAi;
output [162:162] b6_2ZTGIf;

    wire b3_P_F_6_bm_46, b3_P_F_6_am_46, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_46), .B(
        b4_nUAi[488]), .C(b3_P_F_6_am_46), .Y(b6_2ZTGIf[162]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[162]), .B(
        b11_OFWNT9L_8tZ[214]), .C(b4_nUAi[487]), .D(b4_nUAi[486]), .Y(
        b3_P_F_6_am_46));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[162]), .B(
        b11_OFWNT9L_8tZ[214]), .C(b4_nUAi[486]), .D(b4_nUAi[487]), .Y(
        b3_P_F_6_bm_46));
    
endmodule


module b8_1LbcQDr1_x_123_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [253:253] mdiclink_reg;
input  [123:123] b11_OFWNT9L_8tZ;
input  [760:759] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[253]), .B(
        b11_OFWNT9L_8tZ[123]), .C(b4_nUAi[760]), .D(b4_nUAi[759]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[253]), .B(
        b11_OFWNT9L_8tZ[123]), .C(b4_nUAi[760]), .D(b4_nUAi[759]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_324_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [52:52] mdiclink_reg;
input  [324:324] b11_OFWNT9L_8tZ;
input  [158:156] b4_nUAi;
output [52:52] b6_2ZTGIf;

    wire b3_P_F_6_bm_188, b3_P_F_6_am_188, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_188), .B(
        b4_nUAi[158]), .C(b3_P_F_6_am_188), .Y(b6_2ZTGIf[52]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[52]), .B(
        b11_OFWNT9L_8tZ[324]), .C(b4_nUAi[157]), .D(b4_nUAi[156]), .Y(
        b3_P_F_6_am_188));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[52]), .B(
        b11_OFWNT9L_8tZ[324]), .C(b4_nUAi[156]), .D(b4_nUAi[157]), .Y(
        b3_P_F_6_bm_188));
    
endmodule


module b8_1LbcQDr1_x_131_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [245:245] mdiclink_reg;
input  [131:131] b11_OFWNT9L_8tZ;
input  [736:735] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[245]), .B(
        b11_OFWNT9L_8tZ[131]), .C(b4_nUAi[736]), .D(b4_nUAi[735]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[245]), .B(
        b11_OFWNT9L_8tZ[131]), .C(b4_nUAi[736]), .D(b4_nUAi[735]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_102_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [274:274] mdiclink_reg;
input  [102:102] b11_OFWNT9L_8tZ;
input  [824:822] b4_nUAi;
output [274:274] b6_2ZTGIf;

    wire b3_P_F_6_bm_96, b3_P_F_6_am_96, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_96), .B(
        b4_nUAi[824]), .C(b3_P_F_6_am_96), .Y(b6_2ZTGIf[274]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[274]), .B(
        b11_OFWNT9L_8tZ[102]), .C(b4_nUAi[823]), .D(b4_nUAi[822]), .Y(
        b3_P_F_6_am_96));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[274]), .B(
        b11_OFWNT9L_8tZ[102]), .C(b4_nUAi[822]), .D(b4_nUAi[823]), .Y(
        b3_P_F_6_bm_96));
    
endmodule


module b8_1LbcQDr1_x_234_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [142:142] mdiclink_reg;
input  [234:234] b11_OFWNT9L_8tZ;
input  [427:426] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[142]), .B(
        b11_OFWNT9L_8tZ[234]), .C(b4_nUAi[427]), .D(b4_nUAi[426]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[142]), .B(
        b11_OFWNT9L_8tZ[234]), .C(b4_nUAi[427]), .D(b4_nUAi[426]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_160_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [216:216] mdiclink_reg;
input  [160:160] b11_OFWNT9L_8tZ;
input  [650:648] b4_nUAi;
output [216:216] b6_2ZTGIf;

    wire b3_P_F_6_bm_71, b3_P_F_6_am_71, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_71), .B(
        b4_nUAi[650]), .C(b3_P_F_6_am_71), .Y(b6_2ZTGIf[216]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[216]), .B(
        b11_OFWNT9L_8tZ[160]), .C(b4_nUAi[649]), .D(b4_nUAi[648]), .Y(
        b3_P_F_6_am_71));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[216]), .B(
        b11_OFWNT9L_8tZ[160]), .C(b4_nUAi[648]), .D(b4_nUAi[649]), .Y(
        b3_P_F_6_bm_71));
    
endmodule


module b8_1LbcQDr1_x_283_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [93:93] mdiclink_reg;
input  [283:283] b11_OFWNT9L_8tZ;
input  [280:279] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[93]), .B(
        b11_OFWNT9L_8tZ[283]), .C(b4_nUAi[280]), .D(b4_nUAi[279]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[93]), .B(
        b11_OFWNT9L_8tZ[283]), .C(b4_nUAi[280]), .D(b4_nUAi[279]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_370_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [6:6] mdiclink_reg;
input  [370:370] b11_OFWNT9L_8tZ;
input  [20:18] b4_nUAi;
output [6:6] b6_2ZTGIf;

    wire b3_P_F_6_bm_157, b3_P_F_6_am_157, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_157), .B(
        b4_nUAi[20]), .C(b3_P_F_6_am_157), .Y(b6_2ZTGIf[6]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[6]), .B(
        b11_OFWNT9L_8tZ[370]), .C(b4_nUAi[19]), .D(b4_nUAi[18]), .Y(
        b3_P_F_6_am_157));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[6]), .B(
        b11_OFWNT9L_8tZ[370]), .C(b4_nUAi[18]), .D(b4_nUAi[19]), .Y(
        b3_P_F_6_bm_157));
    
endmodule


module b8_1LbcQDr1_x_170_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [206:206] mdiclink_reg;
input  [170:170] b11_OFWNT9L_8tZ;
input  [619:618] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[206]), .B(
        b11_OFWNT9L_8tZ[170]), .C(b4_nUAi[619]), .D(b4_nUAi[618]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[206]), .B(
        b11_OFWNT9L_8tZ[170]), .C(b4_nUAi[619]), .D(b4_nUAi[618]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_55_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [321:321] mdiclink_reg;
input  [55:55] b11_OFWNT9L_8tZ;
input  [965:963] b4_nUAi;
output [321:321] b6_2ZTGIf;

    wire b3_P_F_6_bm_127, b3_P_F_6_am_127, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_127), .B(
        b4_nUAi[965]), .C(b3_P_F_6_am_127), .Y(b6_2ZTGIf[321]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[321]), .B(
        b11_OFWNT9L_8tZ[55]), .C(b4_nUAi[964]), .D(b4_nUAi[963]), .Y(
        b3_P_F_6_am_127));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[321]), .B(
        b11_OFWNT9L_8tZ[55]), .C(b4_nUAi[963]), .D(b4_nUAi[964]), .Y(
        b3_P_F_6_bm_127));
    
endmodule


module b8_1LbcQDr1_x_0_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [376:376] mdiclink_reg;
input  [0:0] b11_OFWNT9L_8tZ;
input  [1129:1128] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[376]), .B(
        b11_OFWNT9L_8tZ[0]), .C(b4_nUAi[1129]), .D(b4_nUAi[1128]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[376]), .B(
        b11_OFWNT9L_8tZ[0]), .C(b4_nUAi[1129]), .D(b4_nUAi[1128]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_211_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [165:165] mdiclink_reg;
input  [211:211] b11_OFWNT9L_8tZ;
input  [496:495] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[165]), .B(
        b11_OFWNT9L_8tZ[211]), .C(b4_nUAi[496]), .D(b4_nUAi[495]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[165]), .B(
        b11_OFWNT9L_8tZ[211]), .C(b4_nUAi[496]), .D(b4_nUAi[495]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_192_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [184:184] mdiclink_reg;
input  [192:192] b11_OFWNT9L_8tZ;
input  [554:552] b4_nUAi;
output [184:184] b6_2ZTGIf;

    wire b3_P_F_6_bm_51, b3_P_F_6_am_51, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_51), .B(
        b4_nUAi[554]), .C(b3_P_F_6_am_51), .Y(b6_2ZTGIf[184]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[184]), .B(
        b11_OFWNT9L_8tZ[192]), .C(b4_nUAi[553]), .D(b4_nUAi[552]), .Y(
        b3_P_F_6_am_51));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[184]), .B(
        b11_OFWNT9L_8tZ[192]), .C(b4_nUAi[552]), .D(b4_nUAi[553]), .Y(
        b3_P_F_6_bm_51));
    
endmodule


module b8_1LbcQDr1_x_118_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [258:258] mdiclink_reg;
input  [118:118] b11_OFWNT9L_8tZ;
input  [776:774] b4_nUAi;
output [258:258] b6_2ZTGIf;

    wire b3_P_F_6_bm_86, b3_P_F_6_am_86, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_86), .B(
        b4_nUAi[776]), .C(b3_P_F_6_am_86), .Y(b6_2ZTGIf[258]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[258]), .B(
        b11_OFWNT9L_8tZ[118]), .C(b4_nUAi[775]), .D(b4_nUAi[774]), .Y(
        b3_P_F_6_am_86));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[258]), .B(
        b11_OFWNT9L_8tZ[118]), .C(b4_nUAi[774]), .D(b4_nUAi[775]), .Y(
        b3_P_F_6_bm_86));
    
endmodule


module b8_1LbcQDr1_x_190_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [186:186] mdiclink_reg;
input  [190:190] b11_OFWNT9L_8tZ;
input  [560:558] b4_nUAi;
output [186:186] b6_2ZTGIf;

    wire b3_P_F_6_bm_49, b3_P_F_6_am_49, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_49), .B(
        b4_nUAi[560]), .C(b3_P_F_6_am_49), .Y(b6_2ZTGIf[186]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[186]), .B(
        b11_OFWNT9L_8tZ[190]), .C(b4_nUAi[559]), .D(b4_nUAi[558]), .Y(
        b3_P_F_6_am_49));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[186]), .B(
        b11_OFWNT9L_8tZ[190]), .C(b4_nUAi[558]), .D(b4_nUAi[559]), .Y(
        b3_P_F_6_bm_49));
    
endmodule


module b8_1LbcQDr1_x_153_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [223:223] mdiclink_reg;
input  [153:153] b11_OFWNT9L_8tZ;
input  [670:669] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[223]), .B(
        b11_OFWNT9L_8tZ[153]), .C(b4_nUAi[670]), .D(b4_nUAi[669]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[223]), .B(
        b11_OFWNT9L_8tZ[153]), .C(b4_nUAi[670]), .D(b4_nUAi[669]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_43_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [333:333] mdiclink_reg;
input  [43:43] b11_OFWNT9L_8tZ;
input  [1000:999] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[333]), .B(
        b11_OFWNT9L_8tZ[43]), .C(b4_nUAi[1000]), .D(b4_nUAi[999]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[333]), .B(
        b11_OFWNT9L_8tZ[43]), .C(b4_nUAi[1000]), .D(b4_nUAi[999]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_231_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [145:145] mdiclink_reg;
input  [231:231] b11_OFWNT9L_8tZ;
input  [437:435] b4_nUAi;
output [145:145] b6_2ZTGIf;

    wire b3_P_F_6_bm_37, b3_P_F_6_am_37, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_37), .B(
        b4_nUAi[437]), .C(b3_P_F_6_am_37), .Y(b6_2ZTGIf[145]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[145]), .B(
        b11_OFWNT9L_8tZ[231]), .C(b4_nUAi[436]), .D(b4_nUAi[435]), .Y(
        b3_P_F_6_am_37));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[145]), .B(
        b11_OFWNT9L_8tZ[231]), .C(b4_nUAi[435]), .D(b4_nUAi[436]), .Y(
        b3_P_F_6_bm_37));
    
endmodule


module b8_1LbcQDr1_x_207_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [169:169] mdiclink_reg;
input  [207:207] b11_OFWNT9L_8tZ;
input  [509:507] b4_nUAi;
output [169:169] b6_2ZTGIf;

    wire b3_P_F_6_bm_40, b3_P_F_6_am_40, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_40), .B(
        b4_nUAi[509]), .C(b3_P_F_6_am_40), .Y(b6_2ZTGIf[169]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[169]), .B(
        b11_OFWNT9L_8tZ[207]), .C(b4_nUAi[508]), .D(b4_nUAi[507]), .Y(
        b3_P_F_6_am_40));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[169]), .B(
        b11_OFWNT9L_8tZ[207]), .C(b4_nUAi[507]), .D(b4_nUAi[508]), .Y(
        b3_P_F_6_bm_40));
    
endmodule


module b8_1LbcQDr1_x_87_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [289:289] mdiclink_reg;
input  [87:87] b11_OFWNT9L_8tZ;
input  [869:867] b4_nUAi;
output [289:289] b6_2ZTGIf;

    wire b3_P_F_6_bm_107, b3_P_F_6_am_107, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_107), .B(
        b4_nUAi[869]), .C(b3_P_F_6_am_107), .Y(b6_2ZTGIf[289]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[289]), .B(
        b11_OFWNT9L_8tZ[87]), .C(b4_nUAi[868]), .D(b4_nUAi[867]), .Y(
        b3_P_F_6_am_107));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[289]), .B(
        b11_OFWNT9L_8tZ[87]), .C(b4_nUAi[867]), .D(b4_nUAi[868]), .Y(
        b3_P_F_6_bm_107));
    
endmodule


module b8_1LbcQDr1_x_331_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [45:45] mdiclink_reg;
input  [331:331] b11_OFWNT9L_8tZ;
input  [136:135] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[45]), .B(
        b11_OFWNT9L_8tZ[331]), .C(b4_nUAi[136]), .D(b4_nUAi[135]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[45]), .B(
        b11_OFWNT9L_8tZ[331]), .C(b4_nUAi[136]), .D(b4_nUAi[135]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_182_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [194:194] mdiclink_reg;
input  [182:182] b11_OFWNT9L_8tZ;
input  [584:582] b4_nUAi;
output [194:194] b6_2ZTGIf;

    wire b3_P_F_6_bm_66, b3_P_F_6_am_66, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_66), .B(
        b4_nUAi[584]), .C(b3_P_F_6_am_66), .Y(b6_2ZTGIf[194]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[194]), .B(
        b11_OFWNT9L_8tZ[182]), .C(b4_nUAi[583]), .D(b4_nUAi[582]), .Y(
        b3_P_F_6_am_66));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[194]), .B(
        b11_OFWNT9L_8tZ[182]), .C(b4_nUAi[582]), .D(b4_nUAi[583]), .Y(
        b3_P_F_6_bm_66));
    
endmodule


module b8_1LbcQDr1_x_208_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [168:168] mdiclink_reg;
input  [208:208] b11_OFWNT9L_8tZ;
input  [506:504] b4_nUAi;
output [168:168] b6_2ZTGIf;

    wire b3_P_F_6_bm_41, b3_P_F_6_am_41, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_41), .B(
        b4_nUAi[506]), .C(b3_P_F_6_am_41), .Y(b6_2ZTGIf[168]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[168]), .B(
        b11_OFWNT9L_8tZ[208]), .C(b4_nUAi[505]), .D(b4_nUAi[504]), .Y(
        b3_P_F_6_am_41));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[168]), .B(
        b11_OFWNT9L_8tZ[208]), .C(b4_nUAi[504]), .D(b4_nUAi[505]), .Y(
        b3_P_F_6_bm_41));
    
endmodule


module b8_1LbcQDr1_x_22_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [354:354] mdiclink_reg;
input  [22:22] b11_OFWNT9L_8tZ;
input  [1064:1062] b4_nUAi;
output [354:354] b6_2ZTGIf;

    wire b3_P_F_6_bm_146, b3_P_F_6_am_146, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_146), .B(
        b4_nUAi[1064]), .C(b3_P_F_6_am_146), .Y(b6_2ZTGIf[354]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[354]), .B(
        b11_OFWNT9L_8tZ[22]), .C(b4_nUAi[1063]), .D(b4_nUAi[1062]), .Y(
        b3_P_F_6_am_146));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[354]), .B(
        b11_OFWNT9L_8tZ[22]), .C(b4_nUAi[1062]), .D(b4_nUAi[1063]), .Y(
        b3_P_F_6_bm_146));
    
endmodule


module b8_1LbcQDr1_x_89_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [287:287] mdiclink_reg;
input  [89:89] b11_OFWNT9L_8tZ;
input  [862:861] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[287]), .B(
        b11_OFWNT9L_8tZ[89]), .C(b4_nUAi[862]), .D(b4_nUAi[861]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[287]), .B(
        b11_OFWNT9L_8tZ[89]), .C(b4_nUAi[862]), .D(b4_nUAi[861]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_180_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [196:196] mdiclink_reg;
input  [180:180] b11_OFWNT9L_8tZ;
input  [590:588] b4_nUAi;
output [196:196] b6_2ZTGIf;

    wire b3_P_F_6_bm_64, b3_P_F_6_am_64, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_64), .B(
        b4_nUAi[590]), .C(b3_P_F_6_am_64), .Y(b6_2ZTGIf[196]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[196]), .B(
        b11_OFWNT9L_8tZ[180]), .C(b4_nUAi[589]), .D(b4_nUAi[588]), .Y(
        b3_P_F_6_am_64));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[196]), .B(
        b11_OFWNT9L_8tZ[180]), .C(b4_nUAi[588]), .D(b4_nUAi[589]), .Y(
        b3_P_F_6_bm_64));
    
endmodule


module b8_1LbcQDr1_x_126_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [250:250] mdiclink_reg;
input  [126:126] b11_OFWNT9L_8tZ;
input  [752:750] b4_nUAi;
output [250:250] b6_2ZTGIf;

    wire b3_P_F_6_bm_223, b3_P_F_6_am_223, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_223), .B(
        b4_nUAi[752]), .C(b3_P_F_6_am_223), .Y(b6_2ZTGIf[250]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[250]), .B(
        b11_OFWNT9L_8tZ[126]), .C(b4_nUAi[751]), .D(b4_nUAi[750]), .Y(
        b3_P_F_6_am_223));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[250]), .B(
        b11_OFWNT9L_8tZ[126]), .C(b4_nUAi[750]), .D(b4_nUAi[751]), .Y(
        b3_P_F_6_bm_223));
    
endmodule


module b8_1LbcQDr1_x_227_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [149:149] mdiclink_reg;
input  [227:227] b11_OFWNT9L_8tZ;
input  [448:447] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[149]), .B(
        b11_OFWNT9L_8tZ[227]), .C(b4_nUAi[448]), .D(b4_nUAi[447]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[149]), .B(
        b11_OFWNT9L_8tZ[227]), .C(b4_nUAi[448]), .D(b4_nUAi[447]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_209_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [167:167] mdiclink_reg;
input  [209:209] b11_OFWNT9L_8tZ;
input  [503:501] b4_nUAi;
output [167:167] b6_2ZTGIf;

    wire b3_P_F_6_bm_42, b3_P_F_6_am_42, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_42), .B(
        b4_nUAi[503]), .C(b3_P_F_6_am_42), .Y(b6_2ZTGIf[167]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[167]), .B(
        b11_OFWNT9L_8tZ[209]), .C(b4_nUAi[502]), .D(b4_nUAi[501]), .Y(
        b3_P_F_6_am_42));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[167]), .B(
        b11_OFWNT9L_8tZ[209]), .C(b4_nUAi[501]), .D(b4_nUAi[502]), .Y(
        b3_P_F_6_bm_42));
    
endmodule


module b8_1LbcQDr1_x_285_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [91:91] mdiclink_reg;
input  [285:285] b11_OFWNT9L_8tZ;
input  [274:273] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[91]), .B(
        b11_OFWNT9L_8tZ[285]), .C(b4_nUAi[274]), .D(b4_nUAi[273]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[91]), .B(
        b11_OFWNT9L_8tZ[285]), .C(b4_nUAi[274]), .D(b4_nUAi[273]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_26_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [350:350] mdiclink_reg;
input  [26:26] b11_OFWNT9L_8tZ;
input  [1051:1050] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[350]), .B(
        b11_OFWNT9L_8tZ[26]), .C(b4_nUAi[1051]), .D(b4_nUAi[1050]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[350]), .B(
        b11_OFWNT9L_8tZ[26]), .C(b4_nUAi[1051]), .D(b4_nUAi[1050]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_371_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [5:5] mdiclink_reg;
input  [371:371] b11_OFWNT9L_8tZ;
input  [16:15] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[5]), .B(
        b11_OFWNT9L_8tZ[371]), .C(b4_nUAi[16]), .D(b4_nUAi[15]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[5]), .B(
        b11_OFWNT9L_8tZ[371]), .C(b4_nUAi[16]), .D(b4_nUAi[15]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_228_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [148:148] mdiclink_reg;
input  [228:228] b11_OFWNT9L_8tZ;
input  [446:444] b4_nUAi;
output [148:148] b6_2ZTGIf;

    wire b3_P_F_6_bm_34, b3_P_F_6_am_34, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_34), .B(
        b4_nUAi[446]), .C(b3_P_F_6_am_34), .Y(b6_2ZTGIf[148]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[148]), .B(
        b11_OFWNT9L_8tZ[228]), .C(b4_nUAi[445]), .D(b4_nUAi[444]), .Y(
        b3_P_F_6_am_34));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[148]), .B(
        b11_OFWNT9L_8tZ[228]), .C(b4_nUAi[444]), .D(b4_nUAi[445]), .Y(
        b3_P_F_6_bm_34));
    
endmodule


module b8_1LbcQDr1_x_77_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [299:299] mdiclink_reg;
input  [77:77] b11_OFWNT9L_8tZ;
input  [898:897] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[299]), .B(
        b11_OFWNT9L_8tZ[77]), .C(b4_nUAi[898]), .D(b4_nUAi[897]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[299]), .B(
        b11_OFWNT9L_8tZ[77]), .C(b4_nUAi[898]), .D(b4_nUAi[897]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_286_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [90:90] mdiclink_reg;
input  [286:286] b11_OFWNT9L_8tZ;
input  [272:270] b4_nUAi;
output [90:90] b6_2ZTGIf;

    wire b3_P_F_6_bm_203, b3_P_F_6_am_203, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_203), .B(
        b4_nUAi[272]), .C(b3_P_F_6_am_203), .Y(b6_2ZTGIf[90]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[90]), .B(
        b11_OFWNT9L_8tZ[286]), .C(b4_nUAi[271]), .D(b4_nUAi[270]), .Y(
        b3_P_F_6_am_203));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[90]), .B(
        b11_OFWNT9L_8tZ[286]), .C(b4_nUAi[270]), .D(b4_nUAi[271]), .Y(
        b3_P_F_6_bm_203));
    
endmodule


module b8_1LbcQDr1_x_141_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [235:235] mdiclink_reg;
input  [141:141] b11_OFWNT9L_8tZ;
input  [706:705] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[235]), .B(
        b11_OFWNT9L_8tZ[141]), .C(b4_nUAi[706]), .D(b4_nUAi[705]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[235]), .B(
        b11_OFWNT9L_8tZ[141]), .C(b4_nUAi[706]), .D(b4_nUAi[705]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_104_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [272:272] mdiclink_reg;
input  [104:104] b11_OFWNT9L_8tZ;
input  [818:816] b4_nUAi;
output [272:272] b6_2ZTGIf;

    wire b3_P_F_6_bm_98, b3_P_F_6_am_98, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_98), .B(
        b4_nUAi[818]), .C(b3_P_F_6_am_98), .Y(b6_2ZTGIf[272]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[272]), .B(
        b11_OFWNT9L_8tZ[104]), .C(b4_nUAi[817]), .D(b4_nUAi[816]), .Y(
        b3_P_F_6_am_98));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[272]), .B(
        b11_OFWNT9L_8tZ[104]), .C(b4_nUAi[816]), .D(b4_nUAi[817]), .Y(
        b3_P_F_6_bm_98));
    
endmodule


module b8_1LbcQDr1_x_216_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [160:160] mdiclink_reg;
input  [216:216] b11_OFWNT9L_8tZ;
input  [482:480] b4_nUAi;
output [160:160] b6_2ZTGIf;

    wire b3_P_F_6_bm_48, b3_P_F_6_am_48, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_48), .B(
        b4_nUAi[482]), .C(b3_P_F_6_am_48), .Y(b6_2ZTGIf[160]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[160]), .B(
        b11_OFWNT9L_8tZ[216]), .C(b4_nUAi[481]), .D(b4_nUAi[480]), .Y(
        b3_P_F_6_am_48));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[160]), .B(
        b11_OFWNT9L_8tZ[216]), .C(b4_nUAi[480]), .D(b4_nUAi[481]), .Y(
        b3_P_F_6_bm_48));
    
endmodule


module b8_1LbcQDr1_x_148_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [228:228] mdiclink_reg;
input  [148:148] b11_OFWNT9L_8tZ;
input  [686:684] b4_nUAi;
output [228:228] b6_2ZTGIf;

    wire b3_P_F_6_bm_218, b3_P_F_6_am_218, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_218), .B(
        b4_nUAi[686]), .C(b3_P_F_6_am_218), .Y(b6_2ZTGIf[228]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[228]), .B(
        b11_OFWNT9L_8tZ[148]), .C(b4_nUAi[685]), .D(b4_nUAi[684]), .Y(
        b3_P_F_6_am_218));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[228]), .B(
        b11_OFWNT9L_8tZ[148]), .C(b4_nUAi[684]), .D(b4_nUAi[685]), .Y(
        b3_P_F_6_bm_218));
    
endmodule


module b8_1LbcQDr1_x_244_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [132:132] mdiclink_reg;
input  [244:244] b11_OFWNT9L_8tZ;
input  [398:396] b4_nUAi;
output [132:132] b6_2ZTGIf;

    wire b3_P_F_6_bm_24, b3_P_F_6_am_24, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_24), .B(
        b4_nUAi[398]), .C(b3_P_F_6_am_24), .Y(b6_2ZTGIf[132]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[132]), .B(
        b11_OFWNT9L_8tZ[244]), .C(b4_nUAi[397]), .D(b4_nUAi[396]), .Y(
        b3_P_F_6_am_24));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[132]), .B(
        b11_OFWNT9L_8tZ[244]), .C(b4_nUAi[396]), .D(b4_nUAi[397]), .Y(
        b3_P_F_6_bm_24));
    
endmodule


module b8_1LbcQDr1_x_79_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [297:297] mdiclink_reg;
input  [79:79] b11_OFWNT9L_8tZ;
input  [893:891] b4_nUAi;
output [297:297] b6_2ZTGIf;

    wire b3_P_F_6_bm_100, b3_P_F_6_am_100, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_100), .B(
        b4_nUAi[893]), .C(b3_P_F_6_am_100), .Y(b6_2ZTGIf[297]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[297]), .B(
        b11_OFWNT9L_8tZ[79]), .C(b4_nUAi[892]), .D(b4_nUAi[891]), .Y(
        b3_P_F_6_am_100));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[297]), .B(
        b11_OFWNT9L_8tZ[79]), .C(b4_nUAi[891]), .D(b4_nUAi[892]), .Y(
        b3_P_F_6_bm_100));
    
endmodule


module b8_1LbcQDr1_x_229_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [147:147] mdiclink_reg;
input  [229:229] b11_OFWNT9L_8tZ;
input  [443:441] b4_nUAi;
output [147:147] b6_2ZTGIf;

    wire b3_P_F_6_bm_35, b3_P_F_6_am_35, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_35), .B(
        b4_nUAi[443]), .C(b3_P_F_6_am_35), .Y(b6_2ZTGIf[147]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[147]), .B(
        b11_OFWNT9L_8tZ[229]), .C(b4_nUAi[442]), .D(b4_nUAi[441]), .Y(
        b3_P_F_6_am_35));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[147]), .B(
        b11_OFWNT9L_8tZ[229]), .C(b4_nUAi[441]), .D(b4_nUAi[442]), .Y(
        b3_P_F_6_bm_35));
    
endmodule


module b8_1LbcQDr1_x_299_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [77:77] mdiclink_reg;
input  [299:299] b11_OFWNT9L_8tZ;
input  [232:231] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[77]), .B(
        b11_OFWNT9L_8tZ[299]), .C(b4_nUAi[232]), .D(b4_nUAi[231]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[77]), .B(
        b11_OFWNT9L_8tZ[299]), .C(b4_nUAi[232]), .D(b4_nUAi[231]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_359_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [17:17] mdiclink_reg;
input  [359:359] b11_OFWNT9L_8tZ;
input  [53:51] b4_nUAi;
output [17:17] b6_2ZTGIf;

    wire b3_P_F_6_bm_171, b3_P_F_6_am_171, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_171), .B(
        b4_nUAi[53]), .C(b3_P_F_6_am_171), .Y(b6_2ZTGIf[17]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[17]), .B(
        b11_OFWNT9L_8tZ[359]), .C(b4_nUAi[52]), .D(b4_nUAi[51]), .Y(
        b3_P_F_6_am_171));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[17]), .B(
        b11_OFWNT9L_8tZ[359]), .C(b4_nUAi[51]), .D(b4_nUAi[52]), .Y(
        b3_P_F_6_bm_171));
    
endmodule


module b8_1LbcQDr1_x_322_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [54:54] mdiclink_reg;
input  [322:322] b11_OFWNT9L_8tZ;
input  [164:162] b4_nUAi;
output [54:54] b6_2ZTGIf;

    wire b3_P_F_6_bm_187, b3_P_F_6_am_187, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_187), .B(
        b4_nUAi[164]), .C(b3_P_F_6_am_187), .Y(b6_2ZTGIf[54]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[54]), .B(
        b11_OFWNT9L_8tZ[322]), .C(b4_nUAi[163]), .D(b4_nUAi[162]), .Y(
        b3_P_F_6_am_187));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[54]), .B(
        b11_OFWNT9L_8tZ[322]), .C(b4_nUAi[162]), .D(b4_nUAi[163]), .Y(
        b3_P_F_6_bm_187));
    
endmodule


module b8_1LbcQDr1_x_374_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [2:2] mdiclink_reg;
input  [374:374] b11_OFWNT9L_8tZ;
input  [8:6] b4_nUAi;
output [2:2] b6_2ZTGIf;

    wire b3_P_F_6_bm_160, b3_P_F_6_am_160, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_160), .B(
        b4_nUAi[8]), .C(b3_P_F_6_am_160), .Y(b6_2ZTGIf[2]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[2]), .B(
        b11_OFWNT9L_8tZ[374]), .C(b4_nUAi[7]), .D(b4_nUAi[6]), .Y(
        b3_P_F_6_am_160));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[2]), .B(
        b11_OFWNT9L_8tZ[374]), .C(b4_nUAi[6]), .D(b4_nUAi[7]), .Y(
        b3_P_F_6_bm_160));
    
endmodule


module b8_1LbcQDr1_x_11_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [365:365] mdiclink_reg;
input  [11:11] b11_OFWNT9L_8tZ;
input  [1096:1095] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[365]), .B(
        b11_OFWNT9L_8tZ[11]), .C(b4_nUAi[1096]), .D(b4_nUAi[1095]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[365]), .B(
        b11_OFWNT9L_8tZ[11]), .C(b4_nUAi[1096]), .D(b4_nUAi[1095]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_319_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [57:57] mdiclink_reg;
input  [319:319] b11_OFWNT9L_8tZ;
input  [173:171] b4_nUAi;
output [57:57] b6_2ZTGIf;

    wire b3_P_F_6_bm_184, b3_P_F_6_am_184, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_184), .B(
        b4_nUAi[173]), .C(b3_P_F_6_am_184), .Y(b6_2ZTGIf[57]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[57]), .B(
        b11_OFWNT9L_8tZ[319]), .C(b4_nUAi[172]), .D(b4_nUAi[171]), .Y(
        b3_P_F_6_am_184));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[57]), .B(
        b11_OFWNT9L_8tZ[319]), .C(b4_nUAi[171]), .D(b4_nUAi[172]), .Y(
        b3_P_F_6_bm_184));
    
endmodule


module b8_1LbcQDr1_x_236_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [140:140] mdiclink_reg;
input  [236:236] b11_OFWNT9L_8tZ;
input  [421:420] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[140]), .B(
        b11_OFWNT9L_8tZ[236]), .C(b4_nUAi[421]), .D(b4_nUAi[420]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[140]), .B(
        b11_OFWNT9L_8tZ[236]), .C(b4_nUAi[421]), .D(b4_nUAi[420]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_338_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [38:38] mdiclink_reg;
input  [338:338] b11_OFWNT9L_8tZ;
input  [116:114] b4_nUAi;
output [38:38] b6_2ZTGIf;

    wire b3_P_F_6_bm_177, b3_P_F_6_am_177, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_177), .B(
        b4_nUAi[116]), .C(b3_P_F_6_am_177), .Y(b6_2ZTGIf[38]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[38]), .B(
        b11_OFWNT9L_8tZ[338]), .C(b4_nUAi[115]), .D(b4_nUAi[114]), .Y(
        b3_P_F_6_am_177));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[38]), .B(
        b11_OFWNT9L_8tZ[338]), .C(b4_nUAi[114]), .D(b4_nUAi[115]), .Y(
        b3_P_F_6_bm_177));
    
endmodule


module b8_1LbcQDr1_x_290_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [86:86] mdiclink_reg;
input  [290:290] b11_OFWNT9L_8tZ;
input  [260:258] b4_nUAi;
output [86:86] b6_2ZTGIf;

    wire b3_P_F_6_bm_207, b3_P_F_6_am_207, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_207), .B(
        b4_nUAi[260]), .C(b3_P_F_6_am_207), .Y(b6_2ZTGIf[86]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[86]), .B(
        b11_OFWNT9L_8tZ[290]), .C(b4_nUAi[259]), .D(b4_nUAi[258]), .Y(
        b3_P_F_6_am_207));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[86]), .B(
        b11_OFWNT9L_8tZ[290]), .C(b4_nUAi[258]), .D(b4_nUAi[259]), .Y(
        b3_P_F_6_bm_207));
    
endmodule


module b8_1LbcQDr1_x_63_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [313:313] mdiclink_reg;
input  [63:63] b11_OFWNT9L_8tZ;
input  [941:939] b4_nUAi;
output [313:313] b6_2ZTGIf;

    wire b3_P_F_6_bm_110, b3_P_F_6_am_110, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_110), .B(
        b4_nUAi[941]), .C(b3_P_F_6_am_110), .Y(b6_2ZTGIf[313]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[313]), .B(
        b11_OFWNT9L_8tZ[63]), .C(b4_nUAi[940]), .D(b4_nUAi[939]), .Y(
        b3_P_F_6_am_110));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[313]), .B(
        b11_OFWNT9L_8tZ[63]), .C(b4_nUAi[939]), .D(b4_nUAi[940]), .Y(
        b3_P_F_6_bm_110));
    
endmodule


module b8_1LbcQDr1_x_334_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [42:42] mdiclink_reg;
input  [334:334] b11_OFWNT9L_8tZ;
input  [128:126] b4_nUAi;
output [42:42] b6_2ZTGIf;

    wire b3_P_F_6_bm_173, b3_P_F_6_am_173, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_173), .B(
        b4_nUAi[128]), .C(b3_P_F_6_am_173), .Y(b6_2ZTGIf[42]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[42]), .B(
        b11_OFWNT9L_8tZ[334]), .C(b4_nUAi[127]), .D(b4_nUAi[126]), .Y(
        b3_P_F_6_am_173));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[42]), .B(
        b11_OFWNT9L_8tZ[334]), .C(b4_nUAi[126]), .D(b4_nUAi[127]), .Y(
        b3_P_F_6_bm_173));
    
endmodule


module b8_1LbcQDr1_x_52_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [324:324] mdiclink_reg;
input  [52:52] b11_OFWNT9L_8tZ;
input  [974:972] b4_nUAi;
output [324:324] b6_2ZTGIf;

    wire b3_P_F_6_bm_124, b3_P_F_6_am_124, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_124), .B(
        b4_nUAi[974]), .C(b3_P_F_6_am_124), .Y(b6_2ZTGIf[324]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[324]), .B(
        b11_OFWNT9L_8tZ[52]), .C(b4_nUAi[973]), .D(b4_nUAi[972]), .Y(
        b3_P_F_6_am_124));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[324]), .B(
        b11_OFWNT9L_8tZ[52]), .C(b4_nUAi[972]), .D(b4_nUAi[973]), .Y(
        b3_P_F_6_bm_124));
    
endmodule


module b8_1LbcQDr1_x_73_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [303:303] mdiclink_reg;
input  [73:73] b11_OFWNT9L_8tZ;
input  [910:909] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[303]), .B(
        b11_OFWNT9L_8tZ[73]), .C(b4_nUAi[910]), .D(b4_nUAi[909]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[303]), .B(
        b11_OFWNT9L_8tZ[73]), .C(b4_nUAi[910]), .D(b4_nUAi[909]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_31_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [345:345] mdiclink_reg;
input  [31:31] b11_OFWNT9L_8tZ;
input  [1037:1035] b4_nUAi;
output [345:345] b6_2ZTGIf;

    wire b3_P_F_6_bm_130, b3_P_F_6_am_130, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_130), .B(
        b4_nUAi[1037]), .C(b3_P_F_6_am_130), .Y(b6_2ZTGIf[345]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[345]), .B(
        b11_OFWNT9L_8tZ[31]), .C(b4_nUAi[1036]), .D(b4_nUAi[1035]), .Y(
        b3_P_F_6_am_130));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[345]), .B(
        b11_OFWNT9L_8tZ[31]), .C(b4_nUAi[1035]), .D(b4_nUAi[1036]), .Y(
        b3_P_F_6_bm_130));
    
endmodule


module b8_1LbcQDr1_x_156_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [220:220] mdiclink_reg;
input  [156:156] b11_OFWNT9L_8tZ;
input  [661:660] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[220]), .B(
        b11_OFWNT9L_8tZ[156]), .C(b4_nUAi[661]), .D(b4_nUAi[660]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[220]), .B(
        b11_OFWNT9L_8tZ[156]), .C(b4_nUAi[661]), .D(b4_nUAi[660]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_215_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [161:161] mdiclink_reg;
input  [215:215] b11_OFWNT9L_8tZ;
input  [485:483] b4_nUAi;
output [161:161] b6_2ZTGIf;

    wire b3_P_F_6_bm_47, b3_P_F_6_am_47, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_47), .B(
        b4_nUAi[485]), .C(b3_P_F_6_am_47), .Y(b6_2ZTGIf[161]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[161]), .B(
        b11_OFWNT9L_8tZ[215]), .C(b4_nUAi[484]), .D(b4_nUAi[483]), .Y(
        b3_P_F_6_am_47));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[161]), .B(
        b11_OFWNT9L_8tZ[215]), .C(b4_nUAi[483]), .D(b4_nUAi[484]), .Y(
        b3_P_F_6_bm_47));
    
endmodule


module b8_1LbcQDr1_x_5_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [371:371] mdiclink_reg;
input  [5:5] b11_OFWNT9L_8tZ;
input  [1115:1113] b4_nUAi;
output [371:371] b6_2ZTGIf;

    wire b3_P_F_6_bm_151, b3_P_F_6_am_151, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_151), .B(
        b4_nUAi[1115]), .C(b3_P_F_6_am_151), .Y(b6_2ZTGIf[371]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[371]), .B(
        b11_OFWNT9L_8tZ[5]), .C(b4_nUAi[1114]), .D(b4_nUAi[1113]), .Y(
        b3_P_F_6_am_151));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[371]), .B(
        b11_OFWNT9L_8tZ[5]), .C(b4_nUAi[1113]), .D(b4_nUAi[1114]), .Y(
        b3_P_F_6_bm_151));
    
endmodule


module b8_1LbcQDr1_x_18_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [358:358] mdiclink_reg;
input  [18:18] b11_OFWNT9L_8tZ;
input  [1076:1074] b4_nUAi;
output [358:358] b6_2ZTGIf;

    wire b3_P_F_6_bm_143, b3_P_F_6_am_143, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_143), .B(
        b4_nUAi[1076]), .C(b3_P_F_6_am_143), .Y(b6_2ZTGIf[358]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[358]), .B(
        b11_OFWNT9L_8tZ[18]), .C(b4_nUAi[1075]), .D(b4_nUAi[1074]), .Y(
        b3_P_F_6_am_143));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[358]), .B(
        b11_OFWNT9L_8tZ[18]), .C(b4_nUAi[1074]), .D(b4_nUAi[1075]), .Y(
        b3_P_F_6_bm_143));
    
endmodule


module b8_1LbcQDr1_x_241_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [135:135] mdiclink_reg;
input  [241:241] b11_OFWNT9L_8tZ;
input  [407:405] b4_nUAi;
output [135:135] b6_2ZTGIf;

    wire b3_P_F_6_bm_22, b3_P_F_6_am_22, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_22), .B(
        b4_nUAi[407]), .C(b3_P_F_6_am_22), .Y(b6_2ZTGIf[135]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[135]), .B(
        b11_OFWNT9L_8tZ[241]), .C(b4_nUAi[406]), .D(b4_nUAi[405]), .Y(
        b3_P_F_6_am_22));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[135]), .B(
        b11_OFWNT9L_8tZ[241]), .C(b4_nUAi[405]), .D(b4_nUAi[406]), .Y(
        b3_P_F_6_bm_22));
    
endmodule


module b8_1LbcQDr1_x_56_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [320:320] mdiclink_reg;
input  [56:56] b11_OFWNT9L_8tZ;
input  [962:960] b4_nUAi;
output [320:320] b6_2ZTGIf;

    wire b3_P_F_6_bm_128, b3_P_F_6_am_128, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_128), .B(
        b4_nUAi[962]), .C(b3_P_F_6_am_128), .Y(b6_2ZTGIf[320]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[320]), .B(
        b11_OFWNT9L_8tZ[56]), .C(b4_nUAi[961]), .D(b4_nUAi[960]), .Y(
        b3_P_F_6_am_128));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[320]), .B(
        b11_OFWNT9L_8tZ[56]), .C(b4_nUAi[960]), .D(b4_nUAi[961]), .Y(
        b3_P_F_6_bm_128));
    
endmodule


module b8_1LbcQDr1_x_14_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [362:362] mdiclink_reg;
input  [14:14] b11_OFWNT9L_8tZ;
input  [1088:1086] b4_nUAi;
output [362:362] b6_2ZTGIf;

    wire b3_P_F_6_bm_139, b3_P_F_6_am_139, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_139), .B(
        b4_nUAi[1088]), .C(b3_P_F_6_am_139), .Y(b6_2ZTGIf[362]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[362]), .B(
        b11_OFWNT9L_8tZ[14]), .C(b4_nUAi[1087]), .D(b4_nUAi[1086]), .Y(
        b3_P_F_6_am_139));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[362]), .B(
        b11_OFWNT9L_8tZ[14]), .C(b4_nUAi[1086]), .D(b4_nUAi[1087]), .Y(
        b3_P_F_6_bm_139));
    
endmodule


module b8_1LbcQDr1_x_337_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [39:39] mdiclink_reg;
input  [337:337] b11_OFWNT9L_8tZ;
input  [119:117] b4_nUAi;
output [39:39] b6_2ZTGIf;

    wire b3_P_F_6_bm_176, b3_P_F_6_am_176, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_176), .B(
        b4_nUAi[119]), .C(b3_P_F_6_am_176), .Y(b6_2ZTGIf[39]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[39]), .B(
        b11_OFWNT9L_8tZ[337]), .C(b4_nUAi[118]), .D(b4_nUAi[117]), .Y(
        b3_P_F_6_am_176));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[39]), .B(
        b11_OFWNT9L_8tZ[337]), .C(b4_nUAi[117]), .D(b4_nUAi[118]), .Y(
        b3_P_F_6_bm_176));
    
endmodule


module b8_1LbcQDr1_x_90_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [286:286] mdiclink_reg;
input  [90:90] b11_OFWNT9L_8tZ;
input  [859:858] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[286]), .B(
        b11_OFWNT9L_8tZ[90]), .C(b4_nUAi[859]), .D(b4_nUAi[858]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[286]), .B(
        b11_OFWNT9L_8tZ[90]), .C(b4_nUAi[859]), .D(b4_nUAi[858]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_235_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [141:141] mdiclink_reg;
input  [235:235] b11_OFWNT9L_8tZ;
input  [424:423] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[141]), .B(
        b11_OFWNT9L_8tZ[235]), .C(b4_nUAi[424]), .D(b4_nUAi[423]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[141]), .B(
        b11_OFWNT9L_8tZ[235]), .C(b4_nUAi[424]), .D(b4_nUAi[423]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_161_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [215:215] mdiclink_reg;
input  [161:161] b11_OFWNT9L_8tZ;
input  [647:645] b4_nUAi;
output [215:215] b6_2ZTGIf;

    wire b3_P_F_6_bm_72, b3_P_F_6_am_72, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_72), .B(
        b4_nUAi[647]), .C(b3_P_F_6_am_72), .Y(b6_2ZTGIf[215]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[215]), .B(
        b11_OFWNT9L_8tZ[161]), .C(b4_nUAi[646]), .D(b4_nUAi[645]), .Y(
        b3_P_F_6_am_72));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[215]), .B(
        b11_OFWNT9L_8tZ[161]), .C(b4_nUAi[645]), .D(b4_nUAi[646]), .Y(
        b3_P_F_6_bm_72));
    
endmodule


module b8_1LbcQDr1_x_103_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [273:273] mdiclink_reg;
input  [103:103] b11_OFWNT9L_8tZ;
input  [821:819] b4_nUAi;
output [273:273] b6_2ZTGIf;

    wire b3_P_F_6_bm_97, b3_P_F_6_am_97, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_97), .B(
        b4_nUAi[821]), .C(b3_P_F_6_am_97), .Y(b6_2ZTGIf[273]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[273]), .B(
        b11_OFWNT9L_8tZ[103]), .C(b4_nUAi[820]), .D(b4_nUAi[819]), .Y(
        b3_P_F_6_am_97));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[273]), .B(
        b11_OFWNT9L_8tZ[103]), .C(b4_nUAi[819]), .D(b4_nUAi[820]), .Y(
        b3_P_F_6_bm_97));
    
endmodule


module b8_1LbcQDr1_x_34_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [342:342] mdiclink_reg;
input  [34:34] b11_OFWNT9L_8tZ;
input  [1028:1026] b4_nUAi;
output [342:342] b6_2ZTGIf;

    wire b3_P_F_6_bm_133, b3_P_F_6_am_133, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_133), .B(
        b4_nUAi[1028]), .C(b3_P_F_6_am_133), .Y(b6_2ZTGIf[342]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[342]), .B(
        b11_OFWNT9L_8tZ[34]), .C(b4_nUAi[1027]), .D(b4_nUAi[1026]), .Y(
        b3_P_F_6_am_133));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[342]), .B(
        b11_OFWNT9L_8tZ[34]), .C(b4_nUAi[1026]), .D(b4_nUAi[1027]), .Y(
        b3_P_F_6_bm_133));
    
endmodule


module b8_1LbcQDr1_x_237_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [139:139] mdiclink_reg;
input  [237:237] b11_OFWNT9L_8tZ;
input  [418:417] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[139]), .B(
        b11_OFWNT9L_8tZ[237]), .C(b4_nUAi[418]), .D(b4_nUAi[417]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[139]), .B(
        b11_OFWNT9L_8tZ[237]), .C(b4_nUAi[418]), .D(b4_nUAi[417]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_264_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [112:112] mdiclink_reg;
input  [264:264] b11_OFWNT9L_8tZ;
input  [338:336] b4_nUAi;
output [112:112] b6_2ZTGIf;

    wire b3_P_F_6_bm_18, b3_P_F_6_am_18, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_18), .B(
        b4_nUAi[338]), .C(b3_P_F_6_am_18), .Y(b6_2ZTGIf[112]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[112]), .B(
        b11_OFWNT9L_8tZ[264]), .C(b4_nUAi[337]), .D(b4_nUAi[336]), .Y(
        b3_P_F_6_am_18));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[112]), .B(
        b11_OFWNT9L_8tZ[264]), .C(b4_nUAi[336]), .D(b4_nUAi[337]), .Y(
        b3_P_F_6_bm_18));
    
endmodule


module b8_1LbcQDr1_x_171_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [205:205] mdiclink_reg;
input  [171:171] b11_OFWNT9L_8tZ;
input  [616:615] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[205]), .B(
        b11_OFWNT9L_8tZ[171]), .C(b4_nUAi[616]), .D(b4_nUAi[615]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[205]), .B(
        b11_OFWNT9L_8tZ[171]), .C(b4_nUAi[616]), .D(b4_nUAi[615]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_80_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [296:296] mdiclink_reg;
input  [80:80] b11_OFWNT9L_8tZ;
input  [890:888] b4_nUAi;
output [296:296] b6_2ZTGIf;

    wire b3_P_F_6_bm_101, b3_P_F_6_am_101, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_101), .B(
        b4_nUAi[890]), .C(b3_P_F_6_am_101), .Y(b6_2ZTGIf[296]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[296]), .B(
        b11_OFWNT9L_8tZ[80]), .C(b4_nUAi[889]), .D(b4_nUAi[888]), .Y(
        b3_P_F_6_am_101));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[296]), .B(
        b11_OFWNT9L_8tZ[80]), .C(b4_nUAi[888]), .D(b4_nUAi[889]), .Y(
        b3_P_F_6_bm_101));
    
endmodule


module b8_1LbcQDr1_x_222_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [154:154] mdiclink_reg;
input  [222:222] b11_OFWNT9L_8tZ;
input  [464:462] b4_nUAi;
output [154:154] b6_2ZTGIf;

    wire b3_P_F_6_bm_29, b3_P_F_6_am_29, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_29), .B(
        b4_nUAi[464]), .C(b3_P_F_6_am_29), .Y(b6_2ZTGIf[154]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[154]), .B(
        b11_OFWNT9L_8tZ[222]), .C(b4_nUAi[463]), .D(b4_nUAi[462]), .Y(
        b3_P_F_6_am_29));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[154]), .B(
        b11_OFWNT9L_8tZ[222]), .C(b4_nUAi[462]), .D(b4_nUAi[463]), .Y(
        b3_P_F_6_bm_29));
    
endmodule


module b8_1LbcQDr1_x_274_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [102:102] mdiclink_reg;
input  [274:274] b11_OFWNT9L_8tZ;
input  [308:306] b4_nUAi;
output [102:102] b6_2ZTGIf;

    wire b3_P_F_6_bm_3, b3_P_F_6_am_3, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_3), .B(
        b4_nUAi[308]), .C(b3_P_F_6_am_3), .Y(b6_2ZTGIf[102]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[102]), .B(
        b11_OFWNT9L_8tZ[274]), .C(b4_nUAi[307]), .D(b4_nUAi[306]), .Y(
        b3_P_F_6_am_3));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[102]), .B(
        b11_OFWNT9L_8tZ[274]), .C(b4_nUAi[306]), .D(b4_nUAi[307]), .Y(
        b3_P_F_6_bm_3));
    
endmodule


module b8_1LbcQDr1_x_238_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [138:138] mdiclink_reg;
input  [238:238] b11_OFWNT9L_8tZ;
input  [416:414] b4_nUAi;
output [138:138] b6_2ZTGIf;

    wire b3_P_F_6_bm_19, b3_P_F_6_am_19, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_19), .B(
        b4_nUAi[416]), .C(b3_P_F_6_am_19), .Y(b6_2ZTGIf[138]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[138]), .B(
        b11_OFWNT9L_8tZ[238]), .C(b4_nUAi[415]), .D(b4_nUAi[414]), .Y(
        b3_P_F_6_am_19));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[138]), .B(
        b11_OFWNT9L_8tZ[238]), .C(b4_nUAi[414]), .D(b4_nUAi[415]), .Y(
        b3_P_F_6_bm_19));
    
endmodule


module b8_1LbcQDr1_x_220_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [156:156] mdiclink_reg;
input  [220:220] b11_OFWNT9L_8tZ;
input  [469:468] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[156]), .B(
        b11_OFWNT9L_8tZ[220]), .C(b4_nUAi[469]), .D(b4_nUAi[468]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[156]), .B(
        b11_OFWNT9L_8tZ[220]), .C(b4_nUAi[469]), .D(b4_nUAi[468]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_239_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [137:137] mdiclink_reg;
input  [239:239] b11_OFWNT9L_8tZ;
input  [413:411] b4_nUAi;
output [137:137] b6_2ZTGIf;

    wire b3_P_F_6_bm_20, b3_P_F_6_am_20, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_20), .B(
        b4_nUAi[413]), .C(b3_P_F_6_am_20), .Y(b6_2ZTGIf[137]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[137]), .B(
        b11_OFWNT9L_8tZ[239]), .C(b4_nUAi[412]), .D(b4_nUAi[411]), .Y(
        b3_P_F_6_am_20));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[137]), .B(
        b11_OFWNT9L_8tZ[239]), .C(b4_nUAi[411]), .D(b4_nUAi[412]), .Y(
        b3_P_F_6_bm_20));
    
endmodule


module b8_1LbcQDr1_x_48_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [328:328] mdiclink_reg;
input  [48:48] b11_OFWNT9L_8tZ;
input  [986:984] b4_nUAi;
output [328:328] b6_2ZTGIf;

    wire b3_P_F_6_bm_121, b3_P_F_6_am_121, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_121), .B(
        b4_nUAi[986]), .C(b3_P_F_6_am_121), .Y(b6_2ZTGIf[328]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[328]), .B(
        b11_OFWNT9L_8tZ[48]), .C(b4_nUAi[985]), .D(b4_nUAi[984]), .Y(
        b3_P_F_6_am_121));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[328]), .B(
        b11_OFWNT9L_8tZ[48]), .C(b4_nUAi[984]), .D(b4_nUAi[985]), .Y(
        b3_P_F_6_bm_121));
    
endmodule


module b8_1LbcQDr1_x_117_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [259:259] mdiclink_reg;
input  [117:117] b11_OFWNT9L_8tZ;
input  [779:777] b4_nUAi;
output [259:259] b6_2ZTGIf;

    wire b3_P_F_6_bm_85, b3_P_F_6_am_85, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_85), .B(
        b4_nUAi[779]), .C(b3_P_F_6_am_85), .Y(b6_2ZTGIf[259]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[259]), .B(
        b11_OFWNT9L_8tZ[117]), .C(b4_nUAi[778]), .D(b4_nUAi[777]), .Y(
        b3_P_F_6_am_85));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[259]), .B(
        b11_OFWNT9L_8tZ[117]), .C(b4_nUAi[777]), .D(b4_nUAi[778]), .Y(
        b3_P_F_6_bm_85));
    
endmodule


module b8_1LbcQDr1_x_7_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [369:369] mdiclink_reg;
input  [7:7] b11_OFWNT9L_8tZ;
input  [1109:1107] b4_nUAi;
output [369:369] b6_2ZTGIf;

    wire b3_P_F_6_bm_152, b3_P_F_6_am_152, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_152), .B(
        b4_nUAi[1109]), .C(b3_P_F_6_am_152), .Y(b6_2ZTGIf[369]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[369]), .B(
        b11_OFWNT9L_8tZ[7]), .C(b4_nUAi[1108]), .D(b4_nUAi[1107]), .Y(
        b3_P_F_6_am_152));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[369]), .B(
        b11_OFWNT9L_8tZ[7]), .C(b4_nUAi[1107]), .D(b4_nUAi[1108]), .Y(
        b3_P_F_6_bm_152));
    
endmodule


module b8_1LbcQDr1_x_350_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [26:26] mdiclink_reg;
input  [350:350] b11_OFWNT9L_8tZ;
input  [80:78] b4_nUAi;
output [26:26] b6_2ZTGIf;

    wire b3_P_F_6_bm_163, b3_P_F_6_am_163, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_163), .B(
        b4_nUAi[80]), .C(b3_P_F_6_am_163), .Y(b6_2ZTGIf[26]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[26]), .B(
        b11_OFWNT9L_8tZ[350]), .C(b4_nUAi[79]), .D(b4_nUAi[78]), .Y(
        b3_P_F_6_am_163));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[26]), .B(
        b11_OFWNT9L_8tZ[350]), .C(b4_nUAi[78]), .D(b4_nUAi[79]), .Y(
        b3_P_F_6_bm_163));
    
endmodule


module b8_1LbcQDr1_x_376_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [0:0] mdiclink_reg;
input  [376:376] b11_OFWNT9L_8tZ;
input  [2:0] b4_nUAi;
output [0:0] b6_2ZTGIf;

    wire b3_P_F_6_bm_162, b3_P_F_6_am_162, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_162), .B(
        b4_nUAi[2]), .C(b3_P_F_6_am_162), .Y(b6_2ZTGIf[0]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[0]), .B(
        b11_OFWNT9L_8tZ[376]), .C(b4_nUAi[1]), .D(b4_nUAi[0]), .Y(
        b3_P_F_6_am_162));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[0]), .B(
        b11_OFWNT9L_8tZ[376]), .C(b4_nUAi[0]), .D(b4_nUAi[1]), .Y(
        b3_P_F_6_bm_162));
    
endmodule


module b8_1LbcQDr1_x_246_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [130:130] mdiclink_reg;
input  [246:246] b11_OFWNT9L_8tZ;
input  [392:390] b4_nUAi;
output [130:130] b6_2ZTGIf;

    wire b3_P_F_6_bm_26, b3_P_F_6_am_26, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_26), .B(
        b4_nUAi[392]), .C(b3_P_F_6_am_26), .Y(b6_2ZTGIf[130]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[130]), .B(
        b11_OFWNT9L_8tZ[246]), .C(b4_nUAi[391]), .D(b4_nUAi[390]), .Y(
        b3_P_F_6_am_26));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[130]), .B(
        b11_OFWNT9L_8tZ[246]), .C(b4_nUAi[390]), .D(b4_nUAi[391]), .Y(
        b3_P_F_6_bm_26));
    
endmodule


module b8_1LbcQDr1_x_310_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [66:66] mdiclink_reg;
input  [310:310] b11_OFWNT9L_8tZ;
input  [200:198] b4_nUAi;
output [66:66] b6_2ZTGIf;

    wire b3_P_F_6_bm_200, b3_P_F_6_am_200, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_200), .B(
        b4_nUAi[200]), .C(b3_P_F_6_am_200), .Y(b6_2ZTGIf[66]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[66]), .B(
        b11_OFWNT9L_8tZ[310]), .C(b4_nUAi[199]), .D(b4_nUAi[198]), .Y(
        b3_P_F_6_am_200));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[66]), .B(
        b11_OFWNT9L_8tZ[310]), .C(b4_nUAi[198]), .D(b4_nUAi[199]), .Y(
        b3_P_F_6_bm_200));
    
endmodule


module b8_1LbcQDr1_x_119_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [257:257] mdiclink_reg;
input  [119:119] b11_OFWNT9L_8tZ;
input  [773:771] b4_nUAi;
output [257:257] b6_2ZTGIf;

    wire b3_P_F_6_bm_87, b3_P_F_6_am_87, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_87), .B(
        b4_nUAi[773]), .C(b3_P_F_6_am_87), .Y(b6_2ZTGIf[257]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[257]), .B(
        b11_OFWNT9L_8tZ[119]), .C(b4_nUAi[772]), .D(b4_nUAi[771]), .Y(
        b3_P_F_6_am_87));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[257]), .B(
        b11_OFWNT9L_8tZ[119]), .C(b4_nUAi[771]), .D(b4_nUAi[772]), .Y(
        b3_P_F_6_bm_87));
    
endmodule


module b8_1LbcQDr1_x_98_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [278:278] mdiclink_reg;
input  [98:98] b11_OFWNT9L_8tZ;
input  [836:834] b4_nUAi;
output [278:278] b6_2ZTGIf;

    wire b3_P_F_6_bm_93, b3_P_F_6_am_93, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_93), .B(
        b4_nUAi[836]), .C(b3_P_F_6_am_93), .Y(b6_2ZTGIf[278]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[278]), .B(
        b11_OFWNT9L_8tZ[98]), .C(b4_nUAi[835]), .D(b4_nUAi[834]), .Y(
        b3_P_F_6_am_93));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[278]), .B(
        b11_OFWNT9L_8tZ[98]), .C(b4_nUAi[834]), .D(b4_nUAi[835]), .Y(
        b3_P_F_6_bm_93));
    
endmodule


module b8_1LbcQDr1_x_261_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [115:115] mdiclink_reg;
input  [261:261] b11_OFWNT9L_8tZ;
input  [347:345] b4_nUAi;
output [115:115] b6_2ZTGIf;

    wire b3_P_F_6_bm_15, b3_P_F_6_am_15, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_15), .B(
        b4_nUAi[347]), .C(b3_P_F_6_am_15), .Y(b6_2ZTGIf[115]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[115]), .B(
        b11_OFWNT9L_8tZ[261]), .C(b4_nUAi[346]), .D(b4_nUAi[345]), .Y(
        b3_P_F_6_am_15));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[115]), .B(
        b11_OFWNT9L_8tZ[261]), .C(b4_nUAi[345]), .D(b4_nUAi[346]), .Y(
        b3_P_F_6_bm_15));
    
endmodule


module b8_1LbcQDr1_x_271_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [105:105] mdiclink_reg;
input  [271:271] b11_OFWNT9L_8tZ;
input  [317:315] b4_nUAi;
output [105:105] b6_2ZTGIf;

    wire b3_P_F_6_bm_0, b3_P_F_6_am_0, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_0), .B(
        b4_nUAi[317]), .C(b3_P_F_6_am_0), .Y(b6_2ZTGIf[105]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[105]), .B(
        b11_OFWNT9L_8tZ[271]), .C(b4_nUAi[316]), .D(b4_nUAi[315]), .Y(
        b3_P_F_6_am_0));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[105]), .B(
        b11_OFWNT9L_8tZ[271]), .C(b4_nUAi[315]), .D(b4_nUAi[316]), .Y(
        b3_P_F_6_bm_0));
    
endmodule


module b8_1LbcQDr1_x_41_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [335:335] mdiclink_reg;
input  [41:41] b11_OFWNT9L_8tZ;
input  [1006:1005] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[335]), .B(
        b11_OFWNT9L_8tZ[41]), .C(b4_nUAi[1006]), .D(b4_nUAi[1005]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[335]), .B(
        b11_OFWNT9L_8tZ[41]), .C(b4_nUAi[1006]), .D(b4_nUAi[1005]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_278_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [98:98] mdiclink_reg;
input  [278:278] b11_OFWNT9L_8tZ;
input  [296:294] b4_nUAi;
output [98:98] b6_2ZTGIf;

    wire b3_P_F_6_bm_6, b3_P_F_6_am_6, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_6), .B(
        b4_nUAi[296]), .C(b3_P_F_6_am_6), .Y(b6_2ZTGIf[98]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[98]), .B(
        b11_OFWNT9L_8tZ[278]), .C(b4_nUAi[295]), .D(b4_nUAi[294]), .Y(
        b3_P_F_6_am_6));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[98]), .B(
        b11_OFWNT9L_8tZ[278]), .C(b4_nUAi[294]), .D(b4_nUAi[295]), .Y(
        b3_P_F_6_bm_6));
    
endmodule


module b8_1LbcQDr1_x_27_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [349:349] mdiclink_reg;
input  [27:27] b11_OFWNT9L_8tZ;
input  [1048:1047] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[349]), .B(
        b11_OFWNT9L_8tZ[27]), .C(b4_nUAi[1048]), .D(b4_nUAi[1047]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[349]), .B(
        b11_OFWNT9L_8tZ[27]), .C(b4_nUAi[1048]), .D(b4_nUAi[1047]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_293_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [83:83] mdiclink_reg;
input  [293:293] b11_OFWNT9L_8tZ;
input  [251:249] b4_nUAi;
output [83:83] b6_2ZTGIf;

    wire b3_P_F_6_bm_209, b3_P_F_6_am_209, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_209), .B(
        b4_nUAi[251]), .C(b3_P_F_6_am_209), .Y(b6_2ZTGIf[83]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[83]), .B(
        b11_OFWNT9L_8tZ[293]), .C(b4_nUAi[250]), .D(b4_nUAi[249]), .Y(
        b3_P_F_6_am_209));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[83]), .B(
        b11_OFWNT9L_8tZ[293]), .C(b4_nUAi[249]), .D(b4_nUAi[250]), .Y(
        b3_P_F_6_bm_209));
    
endmodule


module b8_1LbcQDr1_x_115_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [261:261] mdiclink_reg;
input  [115:115] b11_OFWNT9L_8tZ;
input  [784:783] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[261]), .B(
        b11_OFWNT9L_8tZ[115]), .C(b4_nUAi[784]), .D(b4_nUAi[783]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[261]), .B(
        b11_OFWNT9L_8tZ[115]), .C(b4_nUAi[784]), .D(b4_nUAi[783]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_252_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [124:124] mdiclink_reg;
input  [252:252] b11_OFWNT9L_8tZ;
input  [373:372] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[124]), .B(
        b11_OFWNT9L_8tZ[252]), .C(b4_nUAi[373]), .D(b4_nUAi[372]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[124]), .B(
        b11_OFWNT9L_8tZ[252]), .C(b4_nUAi[373]), .D(b4_nUAi[372]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_329_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [47:47] mdiclink_reg;
input  [329:329] b11_OFWNT9L_8tZ;
input  [142:141] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[47]), .B(
        b11_OFWNT9L_8tZ[329]), .C(b4_nUAi[142]), .D(b4_nUAi[141]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[47]), .B(
        b11_OFWNT9L_8tZ[329]), .C(b4_nUAi[142]), .D(b4_nUAi[141]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_257_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [119:119] mdiclink_reg;
input  [257:257] b11_OFWNT9L_8tZ;
input  [359:357] b4_nUAi;
output [119:119] b6_2ZTGIf;

    wire b3_P_F_6_bm_12, b3_P_F_6_am_12, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_12), .B(
        b4_nUAi[359]), .C(b3_P_F_6_am_12), .Y(b6_2ZTGIf[119]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[119]), .B(
        b11_OFWNT9L_8tZ[257]), .C(b4_nUAi[358]), .D(b4_nUAi[357]), .Y(
        b3_P_F_6_am_12));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[119]), .B(
        b11_OFWNT9L_8tZ[257]), .C(b4_nUAi[357]), .D(b4_nUAi[358]), .Y(
        b3_P_F_6_bm_12));
    
endmodule


module b8_1LbcQDr1_x_250_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [126:126] mdiclink_reg;
input  [250:250] b11_OFWNT9L_8tZ;
input  [379:378] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[126]), .B(
        b11_OFWNT9L_8tZ[250]), .C(b4_nUAi[379]), .D(b4_nUAi[378]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[126]), .B(
        b11_OFWNT9L_8tZ[250]), .C(b4_nUAi[379]), .D(b4_nUAi[378]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_2_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [374:374] mdiclink_reg;
input  [2:2] b11_OFWNT9L_8tZ;
input  [1123:1122] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[374]), .B(
        b11_OFWNT9L_8tZ[2]), .C(b4_nUAi[1123]), .D(b4_nUAi[1122]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[374]), .B(
        b11_OFWNT9L_8tZ[2]), .C(b4_nUAi[1123]), .D(b4_nUAi[1122]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_245_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [131:131] mdiclink_reg;
input  [245:245] b11_OFWNT9L_8tZ;
input  [395:393] b4_nUAi;
output [131:131] b6_2ZTGIf;

    wire b3_P_F_6_bm_25, b3_P_F_6_am_25, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_25), .B(
        b4_nUAi[395]), .C(b3_P_F_6_am_25), .Y(b6_2ZTGIf[131]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[131]), .B(
        b11_OFWNT9L_8tZ[245]), .C(b4_nUAi[394]), .D(b4_nUAi[393]), .Y(
        b3_P_F_6_am_25));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[131]), .B(
        b11_OFWNT9L_8tZ[245]), .C(b4_nUAi[393]), .D(b4_nUAi[394]), .Y(
        b3_P_F_6_bm_25));
    
endmodule


module b8_1LbcQDr1_x_267_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [109:109] mdiclink_reg;
input  [267:267] b11_OFWNT9L_8tZ;
input  [328:327] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[109]), .B(
        b11_OFWNT9L_8tZ[267]), .C(b4_nUAi[328]), .D(b4_nUAi[327]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[109]), .B(
        b11_OFWNT9L_8tZ[267]), .C(b4_nUAi[328]), .D(b4_nUAi[327]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_106_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [270:270] mdiclink_reg;
input  [106:106] b11_OFWNT9L_8tZ;
input  [811:810] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[270]), .B(
        b11_OFWNT9L_8tZ[106]), .C(b4_nUAi[811]), .D(b4_nUAi[810]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[270]), .B(
        b11_OFWNT9L_8tZ[106]), .C(b4_nUAi[811]), .D(b4_nUAi[810]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_213_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [163:163] mdiclink_reg;
input  [213:213] b11_OFWNT9L_8tZ;
input  [491:489] b4_nUAi;
output [163:163] b6_2ZTGIf;

    wire b3_P_F_6_bm_45, b3_P_F_6_am_45, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_45), .B(
        b4_nUAi[491]), .C(b3_P_F_6_am_45), .Y(b6_2ZTGIf[163]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[163]), .B(
        b11_OFWNT9L_8tZ[213]), .C(b4_nUAi[490]), .D(b4_nUAi[489]), .Y(
        b3_P_F_6_am_45));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[163]), .B(
        b11_OFWNT9L_8tZ[213]), .C(b4_nUAi[489]), .D(b4_nUAi[490]), .Y(
        b3_P_F_6_bm_45));
    
endmodule


module b8_1LbcQDr1_x_135_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [241:241] mdiclink_reg;
input  [135:135] b11_OFWNT9L_8tZ;
input  [725:723] b4_nUAi;
output [241:241] b6_2ZTGIf;

    wire b3_P_F_6_bm_231, b3_P_F_6_am_231, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_231), .B(
        b4_nUAi[725]), .C(b3_P_F_6_am_231), .Y(b6_2ZTGIf[241]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[241]), .B(
        b11_OFWNT9L_8tZ[135]), .C(b4_nUAi[724]), .D(b4_nUAi[723]), .Y(
        b3_P_F_6_am_231));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[241]), .B(
        b11_OFWNT9L_8tZ[135]), .C(b4_nUAi[723]), .D(b4_nUAi[724]), .Y(
        b3_P_F_6_bm_231));
    
endmodule


module b8_1LbcQDr1_x_258_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [118:118] mdiclink_reg;
input  [258:258] b11_OFWNT9L_8tZ;
input  [356:354] b4_nUAi;
output [118:118] b6_2ZTGIf;

    wire b3_P_F_6_bm_13, b3_P_F_6_am_13, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_13), .B(
        b4_nUAi[356]), .C(b3_P_F_6_am_13), .Y(b6_2ZTGIf[118]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[118]), .B(
        b11_OFWNT9L_8tZ[258]), .C(b4_nUAi[355]), .D(b4_nUAi[354]), .Y(
        b3_P_F_6_am_13));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[118]), .B(
        b11_OFWNT9L_8tZ[258]), .C(b4_nUAi[354]), .D(b4_nUAi[355]), .Y(
        b3_P_F_6_bm_13));
    
endmodule


module b8_1LbcQDr1_x_277_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [99:99] mdiclink_reg;
input  [277:277] b11_OFWNT9L_8tZ;
input  [299:297] b4_nUAi;
output [99:99] b6_2ZTGIf;

    wire b3_P_F_6_bm_5, b3_P_F_6_am_5, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_5), .B(
        b4_nUAi[299]), .C(b3_P_F_6_am_5), .Y(b6_2ZTGIf[99]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[99]), .B(
        b11_OFWNT9L_8tZ[277]), .C(b4_nUAi[298]), .D(b4_nUAi[297]), .Y(
        b3_P_F_6_am_5));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[99]), .B(
        b11_OFWNT9L_8tZ[277]), .C(b4_nUAi[297]), .D(b4_nUAi[298]), .Y(
        b3_P_F_6_bm_5));
    
endmodule


module b8_1LbcQDr1_x_44_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [332:332] mdiclink_reg;
input  [44:44] b11_OFWNT9L_8tZ;
input  [997:996] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[332]), .B(
        b11_OFWNT9L_8tZ[44]), .C(b4_nUAi[997]), .D(b4_nUAi[996]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[332]), .B(
        b11_OFWNT9L_8tZ[44]), .C(b4_nUAi[997]), .D(b4_nUAi[996]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_341_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [35:35] mdiclink_reg;
input  [341:341] b11_OFWNT9L_8tZ;
input  [107:105] b4_nUAi;
output [35:35] b6_2ZTGIf;

    wire b3_P_F_6_bm_179, b3_P_F_6_am_179, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_179), .B(
        b4_nUAi[107]), .C(b3_P_F_6_am_179), .Y(b6_2ZTGIf[35]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[35]), .B(
        b11_OFWNT9L_8tZ[341]), .C(b4_nUAi[106]), .D(b4_nUAi[105]), .Y(
        b3_P_F_6_am_179));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[35]), .B(
        b11_OFWNT9L_8tZ[341]), .C(b4_nUAi[105]), .D(b4_nUAi[106]), .Y(
        b3_P_F_6_bm_179));
    
endmodule


module b8_1LbcQDr1_x_147_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [229:229] mdiclink_reg;
input  [147:147] b11_OFWNT9L_8tZ;
input  [688:687] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[229]), .B(
        b11_OFWNT9L_8tZ[147]), .C(b4_nUAi[688]), .D(b4_nUAi[687]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[229]), .B(
        b11_OFWNT9L_8tZ[147]), .C(b4_nUAi[688]), .D(b4_nUAi[687]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_268_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [108:108] mdiclink_reg;
input  [268:268] b11_OFWNT9L_8tZ;
input  [325:324] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[108]), .B(
        b11_OFWNT9L_8tZ[268]), .C(b4_nUAi[325]), .D(b4_nUAi[324]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[108]), .B(
        b11_OFWNT9L_8tZ[268]), .C(b4_nUAi[325]), .D(b4_nUAi[324]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_6_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [370:370] mdiclink_reg;
input  [6:6] b11_OFWNT9L_8tZ;
input  [1111:1110] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[370]), .B(
        b11_OFWNT9L_8tZ[6]), .C(b4_nUAi[1111]), .D(b4_nUAi[1110]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[370]), .B(
        b11_OFWNT9L_8tZ[6]), .C(b4_nUAi[1111]), .D(b4_nUAi[1110]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_373_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [3:3] mdiclink_reg;
input  [373:373] b11_OFWNT9L_8tZ;
input  [11:9] b4_nUAi;
output [3:3] b6_2ZTGIf;

    wire b3_P_F_6_bm_159, b3_P_F_6_am_159, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_159), .B(
        b4_nUAi[11]), .C(b3_P_F_6_am_159), .Y(b6_2ZTGIf[3]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[3]), .B(
        b11_OFWNT9L_8tZ[373]), .C(b4_nUAi[10]), .D(b4_nUAi[9]), .Y(
        b3_P_F_6_am_159));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[3]), .B(
        b11_OFWNT9L_8tZ[373]), .C(b4_nUAi[9]), .D(b4_nUAi[10]), .Y(
        b3_P_F_6_bm_159));
    
endmodule


module b8_1LbcQDr1_x_259_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [117:117] mdiclink_reg;
input  [259:259] b11_OFWNT9L_8tZ;
input  [352:351] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[117]), .B(
        b11_OFWNT9L_8tZ[259]), .C(b4_nUAi[352]), .D(b4_nUAi[351]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[117]), .B(
        b11_OFWNT9L_8tZ[259]), .C(b4_nUAi[352]), .D(b4_nUAi[351]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_149_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [227:227] mdiclink_reg;
input  [149:149] b11_OFWNT9L_8tZ;
input  [683:681] b4_nUAi;
output [227:227] b6_2ZTGIf;

    wire b3_P_F_6_bm_219, b3_P_F_6_am_219, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_219), .B(
        b4_nUAi[683]), .C(b3_P_F_6_am_219), .Y(b6_2ZTGIf[227]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[227]), .B(
        b11_OFWNT9L_8tZ[149]), .C(b4_nUAi[682]), .D(b4_nUAi[681]), .Y(
        b3_P_F_6_am_219));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[227]), .B(
        b11_OFWNT9L_8tZ[149]), .C(b4_nUAi[681]), .D(b4_nUAi[682]), .Y(
        b3_P_F_6_bm_219));
    
endmodule


module b8_1LbcQDr1_x_233_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [143:143] mdiclink_reg;
input  [233:233] b11_OFWNT9L_8tZ;
input  [430:429] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[143]), .B(
        b11_OFWNT9L_8tZ[233]), .C(b4_nUAi[430]), .D(b4_nUAi[429]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[143]), .B(
        b11_OFWNT9L_8tZ[233]), .C(b4_nUAi[430]), .D(b4_nUAi[429]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_269_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [107:107] mdiclink_reg;
input  [269:269] b11_OFWNT9L_8tZ;
input  [322:321] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[107]), .B(
        b11_OFWNT9L_8tZ[269]), .C(b4_nUAi[322]), .D(b4_nUAi[321]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[107]), .B(
        b11_OFWNT9L_8tZ[269]), .C(b4_nUAi[322]), .D(b4_nUAi[321]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_266_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [110:110] mdiclink_reg;
input  [266:266] b11_OFWNT9L_8tZ;
input  [331:330] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[110]), .B(
        b11_OFWNT9L_8tZ[266]), .C(b4_nUAi[331]), .D(b4_nUAi[330]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[110]), .B(
        b11_OFWNT9L_8tZ[266]), .C(b4_nUAi[331]), .D(b4_nUAi[330]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_276_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [100:100] mdiclink_reg;
input  [276:276] b11_OFWNT9L_8tZ;
input  [302:300] b4_nUAi;
output [100:100] b6_2ZTGIf;

    wire b3_P_F_6_bm_4, b3_P_F_6_am_4, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_4), .B(
        b4_nUAi[302]), .C(b3_P_F_6_am_4), .Y(b6_2ZTGIf[100]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[100]), .B(
        b11_OFWNT9L_8tZ[276]), .C(b4_nUAi[301]), .D(b4_nUAi[300]), .Y(
        b3_P_F_6_am_4));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[100]), .B(
        b11_OFWNT9L_8tZ[276]), .C(b4_nUAi[300]), .D(b4_nUAi[301]), .Y(
        b3_P_F_6_bm_4));
    
endmodule


module b8_1LbcQDr1_x_120_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [256:256] mdiclink_reg;
input  [120:120] b11_OFWNT9L_8tZ;
input  [770:768] b4_nUAi;
output [256:256] b6_2ZTGIf;

    wire b3_P_F_6_bm_88, b3_P_F_6_am_88, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_88), .B(
        b4_nUAi[770]), .C(b3_P_F_6_am_88), .Y(b6_2ZTGIf[256]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[256]), .B(
        b11_OFWNT9L_8tZ[120]), .C(b4_nUAi[769]), .D(b4_nUAi[768]), .Y(
        b3_P_F_6_am_88));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[256]), .B(
        b11_OFWNT9L_8tZ[120]), .C(b4_nUAi[768]), .D(b4_nUAi[769]), .Y(
        b3_P_F_6_bm_88));
    
endmodule


module b8_1LbcQDr1_x_61_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [315:315] mdiclink_reg;
input  [61:61] b11_OFWNT9L_8tZ;
input  [946:945] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[315]), .B(
        b11_OFWNT9L_8tZ[61]), .C(b4_nUAi[946]), .D(b4_nUAi[945]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[315]), .B(
        b11_OFWNT9L_8tZ[61]), .C(b4_nUAi[946]), .D(b4_nUAi[945]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_295_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [81:81] mdiclink_reg;
input  [295:295] b11_OFWNT9L_8tZ;
input  [245:243] b4_nUAi;
output [81:81] b6_2ZTGIf;

    wire b3_P_F_6_bm_211, b3_P_F_6_am_211, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_211), .B(
        b4_nUAi[245]), .C(b3_P_F_6_am_211), .Y(b6_2ZTGIf[81]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[81]), .B(
        b11_OFWNT9L_8tZ[295]), .C(b4_nUAi[244]), .D(b4_nUAi[243]), .Y(
        b3_P_F_6_am_211));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[81]), .B(
        b11_OFWNT9L_8tZ[295]), .C(b4_nUAi[243]), .D(b4_nUAi[244]), .Y(
        b3_P_F_6_bm_211));
    
endmodule


module b8_1LbcQDr1_x_71_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [305:305] mdiclink_reg;
input  [71:71] b11_OFWNT9L_8tZ;
input  [917:915] b4_nUAi;
output [305:305] b6_2ZTGIf;

    wire b3_P_F_6_bm_117, b3_P_F_6_am_117, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_117), .B(
        b4_nUAi[917]), .C(b3_P_F_6_am_117), .Y(b6_2ZTGIf[305]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[305]), .B(
        b11_OFWNT9L_8tZ[71]), .C(b4_nUAi[916]), .D(b4_nUAi[915]), .Y(
        b3_P_F_6_am_117));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[305]), .B(
        b11_OFWNT9L_8tZ[71]), .C(b4_nUAi[915]), .D(b4_nUAi[916]), .Y(
        b3_P_F_6_bm_117));
    
endmodule


module b8_1LbcQDr1_x_91_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [285:285] mdiclink_reg;
input  [91:91] b11_OFWNT9L_8tZ;
input  [856:855] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[285]), .B(
        b11_OFWNT9L_8tZ[91]), .C(b4_nUAi[856]), .D(b4_nUAi[855]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[285]), .B(
        b11_OFWNT9L_8tZ[91]), .C(b4_nUAi[856]), .D(b4_nUAi[855]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_296_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [80:80] mdiclink_reg;
input  [296:296] b11_OFWNT9L_8tZ;
input  [242:240] b4_nUAi;
output [80:80] b6_2ZTGIf;

    wire b3_P_F_6_bm_212, b3_P_F_6_am_212, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_212), .B(
        b4_nUAi[242]), .C(b3_P_F_6_am_212), .Y(b6_2ZTGIf[80]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[80]), .B(
        b11_OFWNT9L_8tZ[296]), .C(b4_nUAi[241]), .D(b4_nUAi[240]), .Y(
        b3_P_F_6_am_212));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[80]), .B(
        b11_OFWNT9L_8tZ[296]), .C(b4_nUAi[240]), .D(b4_nUAi[241]), .Y(
        b3_P_F_6_bm_212));
    
endmodule


module b8_1LbcQDr1_x_194_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [182:182] mdiclink_reg;
input  [194:194] b11_OFWNT9L_8tZ;
input  [548:546] b4_nUAi;
output [182:182] b6_2ZTGIf;

    wire b3_P_F_6_bm_53, b3_P_F_6_am_53, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_53), .B(
        b4_nUAi[548]), .C(b3_P_F_6_am_53), .Y(b6_2ZTGIf[182]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[182]), .B(
        b11_OFWNT9L_8tZ[194]), .C(b4_nUAi[547]), .D(b4_nUAi[546]), .Y(
        b3_P_F_6_am_53));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[182]), .B(
        b11_OFWNT9L_8tZ[194]), .C(b4_nUAi[546]), .D(b4_nUAi[547]), .Y(
        b3_P_F_6_bm_53));
    
endmodule


module b8_1LbcQDr1_x_344_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [32:32] mdiclink_reg;
input  [344:344] b11_OFWNT9L_8tZ;
input  [98:96] b4_nUAi;
output [32:32] b6_2ZTGIf;

    wire b3_P_F_6_bm_182, b3_P_F_6_am_182, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_182), .B(
        b4_nUAi[98]), .C(b3_P_F_6_am_182), .Y(b6_2ZTGIf[32]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[32]), .B(
        b11_OFWNT9L_8tZ[344]), .C(b4_nUAi[97]), .D(b4_nUAi[96]), .Y(
        b3_P_F_6_am_182));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[32]), .B(
        b11_OFWNT9L_8tZ[344]), .C(b4_nUAi[96]), .D(b4_nUAi[97]), .Y(
        b3_P_F_6_bm_182));
    
endmodule


module b8_1LbcQDr1_x_265_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [111:111] mdiclink_reg;
input  [265:265] b11_OFWNT9L_8tZ;
input  [334:333] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[111]), .B(
        b11_OFWNT9L_8tZ[265]), .C(b4_nUAi[334]), .D(b4_nUAi[333]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[111]), .B(
        b11_OFWNT9L_8tZ[265]), .C(b4_nUAi[334]), .D(b4_nUAi[333]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_37_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [339:339] mdiclink_reg;
input  [37:37] b11_OFWNT9L_8tZ;
input  [1019:1017] b4_nUAi;
output [339:339] b6_2ZTGIf;

    wire b3_P_F_6_bm_135, b3_P_F_6_am_135, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_135), .B(
        b4_nUAi[1019]), .C(b3_P_F_6_am_135), .Y(b6_2ZTGIf[339]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[339]), .B(
        b11_OFWNT9L_8tZ[37]), .C(b4_nUAi[1018]), .D(b4_nUAi[1017]), .Y(
        b3_P_F_6_am_135));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[339]), .B(
        b11_OFWNT9L_8tZ[37]), .C(b4_nUAi[1017]), .D(b4_nUAi[1018]), .Y(
        b3_P_F_6_bm_135));
    
endmodule


module b8_1LbcQDr1_x_353_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [23:23] mdiclink_reg;
input  [353:353] b11_OFWNT9L_8tZ;
input  [71:69] b4_nUAi;
output [23:23] b6_2ZTGIf;

    wire b3_P_F_6_bm_166, b3_P_F_6_am_166, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_166), .B(
        b4_nUAi[71]), .C(b3_P_F_6_am_166), .Y(b6_2ZTGIf[23]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[23]), .B(
        b11_OFWNT9L_8tZ[353]), .C(b4_nUAi[70]), .D(b4_nUAi[69]), .Y(
        b3_P_F_6_am_166));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[23]), .B(
        b11_OFWNT9L_8tZ[353]), .C(b4_nUAi[69]), .D(b4_nUAi[70]), .Y(
        b3_P_F_6_bm_166));
    
endmodule


module b8_1LbcQDr1_x_313_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [63:63] mdiclink_reg;
input  [313:313] b11_OFWNT9L_8tZ;
input  [190:189] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[63]), .B(
        b11_OFWNT9L_8tZ[313]), .C(b4_nUAi[190]), .D(b4_nUAi[189]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[63]), .B(
        b11_OFWNT9L_8tZ[313]), .C(b4_nUAi[190]), .D(b4_nUAi[189]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_275_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [101:101] mdiclink_reg;
input  [275:275] b11_OFWNT9L_8tZ;
input  [304:303] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[101]), .B(
        b11_OFWNT9L_8tZ[275]), .C(b4_nUAi[304]), .D(b4_nUAi[303]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[101]), .B(
        b11_OFWNT9L_8tZ[275]), .C(b4_nUAi[304]), .D(b4_nUAi[303]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_64_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [312:312] mdiclink_reg;
input  [64:64] b11_OFWNT9L_8tZ;
input  [938:936] b4_nUAi;
output [312:312] b6_2ZTGIf;

    wire b3_P_F_6_bm_111, b3_P_F_6_am_111, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_111), .B(
        b4_nUAi[938]), .C(b3_P_F_6_am_111), .Y(b6_2ZTGIf[312]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[312]), .B(
        b11_OFWNT9L_8tZ[64]), .C(b4_nUAi[937]), .D(b4_nUAi[936]), .Y(
        b3_P_F_6_am_111));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[312]), .B(
        b11_OFWNT9L_8tZ[64]), .C(b4_nUAi[936]), .D(b4_nUAi[937]), .Y(
        b3_P_F_6_bm_111));
    
endmodule


module b8_1LbcQDr1_x_81_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [295:295] mdiclink_reg;
input  [81:81] b11_OFWNT9L_8tZ;
input  [887:885] b4_nUAi;
output [295:295] b6_2ZTGIf;

    wire b3_P_F_6_bm_102, b3_P_F_6_am_102, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_102), .B(
        b4_nUAi[887]), .C(b3_P_F_6_am_102), .Y(b6_2ZTGIf[295]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[295]), .B(
        b11_OFWNT9L_8tZ[81]), .C(b4_nUAi[886]), .D(b4_nUAi[885]), .Y(
        b3_P_F_6_am_102));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[295]), .B(
        b11_OFWNT9L_8tZ[81]), .C(b4_nUAi[885]), .D(b4_nUAi[886]), .Y(
        b3_P_F_6_bm_102));
    
endmodule


module b8_1LbcQDr1_x_112_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [264:264] mdiclink_reg;
input  [112:112] b11_OFWNT9L_8tZ;
input  [794:792] b4_nUAi;
output [264:264] b6_2ZTGIf;

    wire b3_P_F_6_bm_81, b3_P_F_6_am_81, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_81), .B(
        b4_nUAi[794]), .C(b3_P_F_6_am_81), .Y(b6_2ZTGIf[264]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[264]), .B(
        b11_OFWNT9L_8tZ[112]), .C(b4_nUAi[793]), .D(b4_nUAi[792]), .Y(
        b3_P_F_6_am_81));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[264]), .B(
        b11_OFWNT9L_8tZ[112]), .C(b4_nUAi[792]), .D(b4_nUAi[793]), .Y(
        b3_P_F_6_bm_81));
    
endmodule


module b8_1LbcQDr1_x_74_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [302:302] mdiclink_reg;
input  [74:74] b11_OFWNT9L_8tZ;
input  [907:906] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[302]), .B(
        b11_OFWNT9L_8tZ[74]), .C(b4_nUAi[907]), .D(b4_nUAi[906]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[302]), .B(
        b11_OFWNT9L_8tZ[74]), .C(b4_nUAi[907]), .D(b4_nUAi[906]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_184_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [192:192] mdiclink_reg;
input  [184:184] b11_OFWNT9L_8tZ;
input  [578:576] b4_nUAi;
output [192:192] b6_2ZTGIf;

    wire b3_P_F_6_bm_68, b3_P_F_6_am_68, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_68), .B(
        b4_nUAi[578]), .C(b3_P_F_6_am_68), .Y(b6_2ZTGIf[192]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[192]), .B(
        b11_OFWNT9L_8tZ[184]), .C(b4_nUAi[577]), .D(b4_nUAi[576]), .Y(
        b3_P_F_6_am_68));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[192]), .B(
        b11_OFWNT9L_8tZ[184]), .C(b4_nUAi[576]), .D(b4_nUAi[577]), .Y(
        b3_P_F_6_bm_68));
    
endmodule


module b8_1LbcQDr1_x_145_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [231:231] mdiclink_reg;
input  [145:145] b11_OFWNT9L_8tZ;
input  [695:693] b4_nUAi;
output [231:231] b6_2ZTGIf;

    wire b3_P_F_6_bm_216, b3_P_F_6_am_216, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_216), .B(
        b4_nUAi[695]), .C(b3_P_F_6_am_216), .Y(b6_2ZTGIf[231]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[231]), .B(
        b11_OFWNT9L_8tZ[145]), .C(b4_nUAi[694]), .D(b4_nUAi[693]), .Y(
        b3_P_F_6_am_216));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[231]), .B(
        b11_OFWNT9L_8tZ[145]), .C(b4_nUAi[693]), .D(b4_nUAi[694]), .Y(
        b3_P_F_6_bm_216));
    
endmodule


module b8_1LbcQDr1_x_150_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [226:226] mdiclink_reg;
input  [150:150] b11_OFWNT9L_8tZ;
input  [680:678] b4_nUAi;
output [226:226] b6_2ZTGIf;

    wire b3_P_F_6_bm_220, b3_P_F_6_am_220, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_220), .B(
        b4_nUAi[680]), .C(b3_P_F_6_am_220), .Y(b6_2ZTGIf[226]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[226]), .B(
        b11_OFWNT9L_8tZ[150]), .C(b4_nUAi[679]), .D(b4_nUAi[678]), .Y(
        b3_P_F_6_am_220));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[226]), .B(
        b11_OFWNT9L_8tZ[150]), .C(b4_nUAi[678]), .D(b4_nUAi[679]), .Y(
        b3_P_F_6_bm_220));
    
endmodule


module b8_1LbcQDr1_x_202_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [174:174] mdiclink_reg;
input  [202:202] b11_OFWNT9L_8tZ;
input  [523:522] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[174]), .B(
        b11_OFWNT9L_8tZ[202]), .C(b4_nUAi[523]), .D(b4_nUAi[522]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[174]), .B(
        b11_OFWNT9L_8tZ[202]), .C(b4_nUAi[523]), .D(b4_nUAi[522]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_132_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [244:244] mdiclink_reg;
input  [132:132] b11_OFWNT9L_8tZ;
input  [734:732] b4_nUAi;
output [244:244] b6_2ZTGIf;

    wire b3_P_F_6_bm_228, b3_P_F_6_am_228, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_228), .B(
        b4_nUAi[734]), .C(b3_P_F_6_am_228), .Y(b6_2ZTGIf[244]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[244]), .B(
        b11_OFWNT9L_8tZ[132]), .C(b4_nUAi[733]), .D(b4_nUAi[732]), .Y(
        b3_P_F_6_am_228));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[244]), .B(
        b11_OFWNT9L_8tZ[132]), .C(b4_nUAi[732]), .D(b4_nUAi[733]), .Y(
        b3_P_F_6_bm_228));
    
endmodule


module b8_1LbcQDr1_x_191_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [185:185] mdiclink_reg;
input  [191:191] b11_OFWNT9L_8tZ;
input  [557:555] b4_nUAi;
output [185:185] b6_2ZTGIf;

    wire b3_P_F_6_bm_50, b3_P_F_6_am_50, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_50), .B(
        b4_nUAi[557]), .C(b3_P_F_6_am_50), .Y(b6_2ZTGIf[185]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[185]), .B(
        b11_OFWNT9L_8tZ[191]), .C(b4_nUAi[556]), .D(b4_nUAi[555]), .Y(
        b3_P_F_6_am_50));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[185]), .B(
        b11_OFWNT9L_8tZ[191]), .C(b4_nUAi[555]), .D(b4_nUAi[556]), .Y(
        b3_P_F_6_bm_50));
    
endmodule


module b8_1LbcQDr1_x_200_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [176:176] mdiclink_reg;
input  [200:200] b11_OFWNT9L_8tZ;
input  [530:528] b4_nUAi;
output [176:176] b6_2ZTGIf;

    wire b3_P_F_6_bm_58, b3_P_F_6_am_58, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_58), .B(
        b4_nUAi[530]), .C(b3_P_F_6_am_58), .Y(b6_2ZTGIf[176]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[176]), .B(
        b11_OFWNT9L_8tZ[200]), .C(b4_nUAi[529]), .D(b4_nUAi[528]), .Y(
        b3_P_F_6_am_58));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[176]), .B(
        b11_OFWNT9L_8tZ[200]), .C(b4_nUAi[528]), .D(b4_nUAi[529]), .Y(
        b3_P_F_6_bm_58));
    
endmodule


module b8_1LbcQDr1_x_10_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [366:366] mdiclink_reg;
input  [10:10] b11_OFWNT9L_8tZ;
input  [1099:1098] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[366]), .B(
        b11_OFWNT9L_8tZ[10]), .C(b4_nUAi[1099]), .D(b4_nUAi[1098]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[366]), .B(
        b11_OFWNT9L_8tZ[10]), .C(b4_nUAi[1099]), .D(b4_nUAi[1098]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_243_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [133:133] mdiclink_reg;
input  [243:243] b11_OFWNT9L_8tZ;
input  [400:399] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[133]), .B(
        b11_OFWNT9L_8tZ[243]), .C(b4_nUAi[400]), .D(b4_nUAi[399]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[133]), .B(
        b11_OFWNT9L_8tZ[243]), .C(b4_nUAi[400]), .D(b4_nUAi[399]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_281_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [95:95] mdiclink_reg;
input  [281:281] b11_OFWNT9L_8tZ;
input  [286:285] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[95]), .B(
        b11_OFWNT9L_8tZ[281]), .C(b4_nUAi[286]), .D(b4_nUAi[285]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[95]), .B(
        b11_OFWNT9L_8tZ[281]), .C(b4_nUAi[286]), .D(b4_nUAi[285]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_368_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [8:8] mdiclink_reg;
input  [368:368] b11_OFWNT9L_8tZ;
input  [26:24] b4_nUAi;
output [8:8] b6_2ZTGIf;

    wire b3_P_F_6_bm_155, b3_P_F_6_am_155, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_155), .B(
        b4_nUAi[26]), .C(b3_P_F_6_am_155), .Y(b6_2ZTGIf[8]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[8]), .B(
        b11_OFWNT9L_8tZ[368]), .C(b4_nUAi[25]), .D(b4_nUAi[24]), .Y(
        b3_P_F_6_am_155));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[8]), .B(
        b11_OFWNT9L_8tZ[368]), .C(b4_nUAi[24]), .D(b4_nUAi[25]), .Y(
        b3_P_F_6_bm_155));
    
endmodule


module b8_1LbcQDr1_x_97_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [279:279] mdiclink_reg;
input  [97:97] b11_OFWNT9L_8tZ;
input  [839:837] b4_nUAi;
output [279:279] b6_2ZTGIf;

    wire b3_P_F_6_bm_92, b3_P_F_6_am_92, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_92), .B(
        b4_nUAi[839]), .C(b3_P_F_6_am_92), .Y(b6_2ZTGIf[279]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[279]), .B(
        b11_OFWNT9L_8tZ[97]), .C(b4_nUAi[838]), .D(b4_nUAi[837]), .Y(
        b3_P_F_6_am_92));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[279]), .B(
        b11_OFWNT9L_8tZ[97]), .C(b4_nUAi[837]), .D(b4_nUAi[838]), .Y(
        b3_P_F_6_bm_92));
    
endmodule


module b8_1LbcQDr1_x_30_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [346:346] mdiclink_reg;
input  [30:30] b11_OFWNT9L_8tZ;
input  [1040:1038] b4_nUAi;
output [346:346] b6_2ZTGIf;

    wire b3_P_F_6_bm_129, b3_P_F_6_am_129, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_129), .B(
        b4_nUAi[1040]), .C(b3_P_F_6_am_129), .Y(b6_2ZTGIf[346]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[346]), .B(
        b11_OFWNT9L_8tZ[30]), .C(b4_nUAi[1039]), .D(b4_nUAi[1038]), .Y(
        b3_P_F_6_am_129));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[346]), .B(
        b11_OFWNT9L_8tZ[30]), .C(b4_nUAi[1038]), .D(b4_nUAi[1039]), .Y(
        b3_P_F_6_bm_129));
    
endmodule


module b8_1LbcQDr1_x_187_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [189:189] mdiclink_reg;
input  [187:187] b11_OFWNT9L_8tZ;
input  [568:567] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[189]), .B(
        b11_OFWNT9L_8tZ[187]), .C(b4_nUAi[568]), .D(b4_nUAi[567]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[189]), .B(
        b11_OFWNT9L_8tZ[187]), .C(b4_nUAi[568]), .D(b4_nUAi[567]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_181_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [195:195] mdiclink_reg;
input  [181:181] b11_OFWNT9L_8tZ;
input  [587:585] b4_nUAi;
output [195:195] b6_2ZTGIf;

    wire b3_P_F_6_bm_65, b3_P_F_6_am_65, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_65), .B(
        b4_nUAi[587]), .C(b3_P_F_6_am_65), .Y(b6_2ZTGIf[195]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[195]), .B(
        b11_OFWNT9L_8tZ[181]), .C(b4_nUAi[586]), .D(b4_nUAi[585]), .Y(
        b3_P_F_6_am_65));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[195]), .B(
        b11_OFWNT9L_8tZ[181]), .C(b4_nUAi[585]), .D(b4_nUAi[586]), .Y(
        b3_P_F_6_bm_65));
    
endmodule


module b8_1LbcQDr1_x_99_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [277:277] mdiclink_reg;
input  [99:99] b11_OFWNT9L_8tZ;
input  [832:831] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[277]), .B(
        b11_OFWNT9L_8tZ[99]), .C(b4_nUAi[832]), .D(b4_nUAi[831]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[277]), .B(
        b11_OFWNT9L_8tZ[99]), .C(b4_nUAi[832]), .D(b4_nUAi[831]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_57_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [319:319] mdiclink_reg;
input  [57:57] b11_OFWNT9L_8tZ;
input  [958:957] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[319]), .B(
        b11_OFWNT9L_8tZ[57]), .C(b4_nUAi[958]), .D(b4_nUAi[957]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[319]), .B(
        b11_OFWNT9L_8tZ[57]), .C(b4_nUAi[958]), .D(b4_nUAi[957]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_355_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [21:21] mdiclink_reg;
input  [355:355] b11_OFWNT9L_8tZ;
input  [64:63] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[21]), .B(
        b11_OFWNT9L_8tZ[355]), .C(b4_nUAi[64]), .D(b4_nUAi[63]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[21]), .B(
        b11_OFWNT9L_8tZ[355]), .C(b4_nUAi[64]), .D(b4_nUAi[63]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_188_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [188:188] mdiclink_reg;
input  [188:188] b11_OFWNT9L_8tZ;
input  [565:564] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[188]), .B(
        b11_OFWNT9L_8tZ[188]), .C(b4_nUAi[565]), .D(b4_nUAi[564]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[188]), .B(
        b11_OFWNT9L_8tZ[188]), .C(b4_nUAi[565]), .D(b4_nUAi[564]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_315_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [61:61] mdiclink_reg;
input  [315:315] b11_OFWNT9L_8tZ;
input  [184:183] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[61]), .B(
        b11_OFWNT9L_8tZ[315]), .C(b4_nUAi[184]), .D(b4_nUAi[183]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[61]), .B(
        b11_OFWNT9L_8tZ[315]), .C(b4_nUAi[184]), .D(b4_nUAi[183]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_67_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [309:309] mdiclink_reg;
input  [67:67] b11_OFWNT9L_8tZ;
input  [928:927] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[309]), .B(
        b11_OFWNT9L_8tZ[67]), .C(b4_nUAi[928]), .D(b4_nUAi[927]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[309]), .B(
        b11_OFWNT9L_8tZ[67]), .C(b4_nUAi[928]), .D(b4_nUAi[927]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_9_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [367:367] mdiclink_reg;
input  [9:9] b11_OFWNT9L_8tZ;
input  [1102:1101] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[367]), .B(
        b11_OFWNT9L_8tZ[9]), .C(b4_nUAi[1102]), .D(b4_nUAi[1101]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[367]), .B(
        b11_OFWNT9L_8tZ[9]), .C(b4_nUAi[1102]), .D(b4_nUAi[1101]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_356_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [20:20] mdiclink_reg;
input  [356:356] b11_OFWNT9L_8tZ;
input  [62:60] b4_nUAi;
output [20:20] b6_2ZTGIf;

    wire b3_P_F_6_bm_168, b3_P_F_6_am_168, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_168), .B(
        b4_nUAi[62]), .C(b3_P_F_6_am_168), .Y(b6_2ZTGIf[20]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[20]), .B(
        b11_OFWNT9L_8tZ[356]), .C(b4_nUAi[61]), .D(b4_nUAi[60]), .Y(
        b3_P_F_6_am_168));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[20]), .B(
        b11_OFWNT9L_8tZ[356]), .C(b4_nUAi[60]), .D(b4_nUAi[61]), .Y(
        b3_P_F_6_bm_168));
    
endmodule


module b8_1LbcQDr1_x_23_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [353:353] mdiclink_reg;
input  [23:23] b11_OFWNT9L_8tZ;
input  [1061:1059] b4_nUAi;
output [353:353] b6_2ZTGIf;

    wire b3_P_F_6_bm_147, b3_P_F_6_am_147, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_147), .B(
        b4_nUAi[1061]), .C(b3_P_F_6_am_147), .Y(b6_2ZTGIf[353]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[353]), .B(
        b11_OFWNT9L_8tZ[23]), .C(b4_nUAi[1060]), .D(b4_nUAi[1059]), .Y(
        b3_P_F_6_am_147));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[353]), .B(
        b11_OFWNT9L_8tZ[23]), .C(b4_nUAi[1059]), .D(b4_nUAi[1060]), .Y(
        b3_P_F_6_bm_147));
    
endmodule


module b8_1LbcQDr1_x_316_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [60:60] mdiclink_reg;
input  [316:316] b11_OFWNT9L_8tZ;
input  [181:180] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[60]), .B(
        b11_OFWNT9L_8tZ[316]), .C(b4_nUAi[181]), .D(b4_nUAi[180]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[60]), .B(
        b11_OFWNT9L_8tZ[316]), .C(b4_nUAi[181]), .D(b4_nUAi[180]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_189_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [187:187] mdiclink_reg;
input  [189:189] b11_OFWNT9L_8tZ;
input  [562:561] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[187]), .B(
        b11_OFWNT9L_8tZ[189]), .C(b4_nUAi[562]), .D(b4_nUAi[561]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[187]), .B(
        b11_OFWNT9L_8tZ[189]), .C(b4_nUAi[562]), .D(b4_nUAi[561]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_177_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [199:199] mdiclink_reg;
input  [177:177] b11_OFWNT9L_8tZ;
input  [599:597] b4_nUAi;
output [199:199] b6_2ZTGIf;

    wire b3_P_F_6_bm_62, b3_P_F_6_am_62, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_62), .B(
        b4_nUAi[599]), .C(b3_P_F_6_am_62), .Y(b6_2ZTGIf[199]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[199]), .B(
        b11_OFWNT9L_8tZ[177]), .C(b4_nUAi[598]), .D(b4_nUAi[597]), .Y(
        b3_P_F_6_am_62));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[199]), .B(
        b11_OFWNT9L_8tZ[177]), .C(b4_nUAi[597]), .D(b4_nUAi[598]), .Y(
        b3_P_F_6_bm_62));
    
endmodule


module b8_1LbcQDr1_x_165_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [211:211] mdiclink_reg;
input  [165:165] b11_OFWNT9L_8tZ;
input  [635:633] b4_nUAi;
output [211:211] b6_2ZTGIf;

    wire b3_P_F_6_bm_75, b3_P_F_6_am_75, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_75), .B(
        b4_nUAi[635]), .C(b3_P_F_6_am_75), .Y(b6_2ZTGIf[211]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[211]), .B(
        b11_OFWNT9L_8tZ[165]), .C(b4_nUAi[634]), .D(b4_nUAi[633]), .Y(
        b3_P_F_6_am_75));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[211]), .B(
        b11_OFWNT9L_8tZ[165]), .C(b4_nUAi[633]), .D(b4_nUAi[634]), .Y(
        b3_P_F_6_bm_75));
    
endmodule


module b8_1LbcQDr1_x_29_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [347:347] mdiclink_reg;
input  [29:29] b11_OFWNT9L_8tZ;
input  [1042:1041] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[347]), .B(
        b11_OFWNT9L_8tZ[29]), .C(b4_nUAi[1042]), .D(b4_nUAi[1041]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[347]), .B(
        b11_OFWNT9L_8tZ[29]), .C(b4_nUAi[1042]), .D(b4_nUAi[1041]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_196_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [180:180] mdiclink_reg;
input  [196:196] b11_OFWNT9L_8tZ;
input  [542:540] b4_nUAi;
output [180:180] b6_2ZTGIf;

    wire b3_P_F_6_bm_54, b3_P_F_6_am_54, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_54), .B(
        b4_nUAi[542]), .C(b3_P_F_6_am_54), .Y(b6_2ZTGIf[180]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[180]), .B(
        b11_OFWNT9L_8tZ[196]), .C(b4_nUAi[541]), .D(b4_nUAi[540]), .Y(
        b3_P_F_6_am_54));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[180]), .B(
        b11_OFWNT9L_8tZ[196]), .C(b4_nUAi[540]), .D(b4_nUAi[541]), .Y(
        b3_P_F_6_bm_54));
    
endmodule


module b8_1LbcQDr1_x_114_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [262:262] mdiclink_reg;
input  [114:114] b11_OFWNT9L_8tZ;
input  [788:786] b4_nUAi;
output [262:262] b6_2ZTGIf;

    wire b3_P_F_6_bm_83, b3_P_F_6_am_83, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_83), .B(
        b4_nUAi[788]), .C(b3_P_F_6_am_83), .Y(b6_2ZTGIf[262]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[262]), .B(
        b11_OFWNT9L_8tZ[114]), .C(b4_nUAi[787]), .D(b4_nUAi[786]), .Y(
        b3_P_F_6_am_83));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[262]), .B(
        b11_OFWNT9L_8tZ[114]), .C(b4_nUAi[786]), .D(b4_nUAi[787]), .Y(
        b3_P_F_6_bm_83));
    
endmodule


module b8_1LbcQDr1_x_178_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [198:198] mdiclink_reg;
input  [178:178] b11_OFWNT9L_8tZ;
input  [596:594] b4_nUAi;
output [198:198] b6_2ZTGIf;

    wire b3_P_F_6_bm_63, b3_P_F_6_am_63, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_63), .B(
        b4_nUAi[596]), .C(b3_P_F_6_am_63), .Y(b6_2ZTGIf[198]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[198]), .B(
        b11_OFWNT9L_8tZ[178]), .C(b4_nUAi[595]), .D(b4_nUAi[594]), .Y(
        b3_P_F_6_am_63));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[198]), .B(
        b11_OFWNT9L_8tZ[178]), .C(b4_nUAi[594]), .D(b4_nUAi[595]), .Y(
        b3_P_F_6_bm_63));
    
endmodule


module b8_1LbcQDr1_x_284_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [92:92] mdiclink_reg;
input  [284:284] b11_OFWNT9L_8tZ;
input  [277:276] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[92]), .B(
        b11_OFWNT9L_8tZ[284]), .C(b4_nUAi[277]), .D(b4_nUAi[276]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[92]), .B(
        b11_OFWNT9L_8tZ[284]), .C(b4_nUAi[277]), .D(b4_nUAi[276]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_175_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [201:201] mdiclink_reg;
input  [175:175] b11_OFWNT9L_8tZ;
input  [605:603] b4_nUAi;
output [201:201] b6_2ZTGIf;

    wire b3_P_F_6_bm_60, b3_P_F_6_am_60, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_60), .B(
        b4_nUAi[605]), .C(b3_P_F_6_am_60), .Y(b6_2ZTGIf[201]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[201]), .B(
        b11_OFWNT9L_8tZ[175]), .C(b4_nUAi[604]), .D(b4_nUAi[603]), .Y(
        b3_P_F_6_am_60));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[201]), .B(
        b11_OFWNT9L_8tZ[175]), .C(b4_nUAi[603]), .D(b4_nUAi[604]), .Y(
        b3_P_F_6_bm_60));
    
endmodule


module b8_1LbcQDr1_x_300_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [76:76] mdiclink_reg;
input  [300:300] b11_OFWNT9L_8tZ;
input  [229:228] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[76]), .B(
        b11_OFWNT9L_8tZ[300]), .C(b4_nUAi[229]), .D(b4_nUAi[228]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[76]), .B(
        b11_OFWNT9L_8tZ[300]), .C(b4_nUAi[229]), .D(b4_nUAi[228]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_360_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [16:16] mdiclink_reg;
input  [360:360] b11_OFWNT9L_8tZ;
input  [50:48] b4_nUAi;
output [16:16] b6_2ZTGIf;

    wire b3_P_F_6_bm_172, b3_P_F_6_am_172, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_172), .B(
        b4_nUAi[50]), .C(b3_P_F_6_am_172), .Y(b6_2ZTGIf[16]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[16]), .B(
        b11_OFWNT9L_8tZ[360]), .C(b4_nUAi[49]), .D(b4_nUAi[48]), .Y(
        b3_P_F_6_am_172));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[16]), .B(
        b11_OFWNT9L_8tZ[360]), .C(b4_nUAi[48]), .D(b4_nUAi[49]), .Y(
        b3_P_F_6_bm_172));
    
endmodule


module b8_1LbcQDr1_x_339_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [37:37] mdiclink_reg;
input  [339:339] b11_OFWNT9L_8tZ;
input  [112:111] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[37]), .B(
        b11_OFWNT9L_8tZ[339]), .C(b4_nUAi[112]), .D(b4_nUAi[111]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[37]), .B(
        b11_OFWNT9L_8tZ[339]), .C(b4_nUAi[112]), .D(b4_nUAi[111]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_179_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [197:197] mdiclink_reg;
input  [179:179] b11_OFWNT9L_8tZ;
input  [592:591] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[197]), .B(
        b11_OFWNT9L_8tZ[179]), .C(b4_nUAi[592]), .D(b4_nUAi[591]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[197]), .B(
        b11_OFWNT9L_8tZ[179]), .C(b4_nUAi[592]), .D(b4_nUAi[591]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_263_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [113:113] mdiclink_reg;
input  [263:263] b11_OFWNT9L_8tZ;
input  [341:339] b4_nUAi;
output [113:113] b6_2ZTGIf;

    wire b3_P_F_6_bm_17, b3_P_F_6_am_17, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_17), .B(
        b4_nUAi[341]), .C(b3_P_F_6_am_17), .Y(b6_2ZTGIf[113]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[113]), .B(
        b11_OFWNT9L_8tZ[263]), .C(b4_nUAi[340]), .D(b4_nUAi[339]), .Y(
        b3_P_F_6_am_17));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[113]), .B(
        b11_OFWNT9L_8tZ[263]), .C(b4_nUAi[339]), .D(b4_nUAi[340]), .Y(
        b3_P_F_6_bm_17));
    
endmodule


module b8_1LbcQDr1_x_288_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [88:88] mdiclink_reg;
input  [288:288] b11_OFWNT9L_8tZ;
input  [266:264] b4_nUAi;
output [88:88] b6_2ZTGIf;

    wire b3_P_F_6_bm_205, b3_P_F_6_am_205, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_205), .B(
        b4_nUAi[266]), .C(b3_P_F_6_am_205), .Y(b6_2ZTGIf[88]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[88]), .B(
        b11_OFWNT9L_8tZ[288]), .C(b4_nUAi[265]), .D(b4_nUAi[264]), .Y(
        b3_P_F_6_am_205));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[88]), .B(
        b11_OFWNT9L_8tZ[288]), .C(b4_nUAi[264]), .D(b4_nUAi[265]), .Y(
        b3_P_F_6_bm_205));
    
endmodule


module b8_1LbcQDr1_x_134_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [242:242] mdiclink_reg;
input  [134:134] b11_OFWNT9L_8tZ;
input  [728:726] b4_nUAi;
output [242:242] b6_2ZTGIf;

    wire b3_P_F_6_bm_230, b3_P_F_6_am_230, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_230), .B(
        b4_nUAi[728]), .C(b3_P_F_6_am_230), .Y(b6_2ZTGIf[242]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[242]), .B(
        b11_OFWNT9L_8tZ[134]), .C(b4_nUAi[727]), .D(b4_nUAi[726]), .Y(
        b3_P_F_6_am_230));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[242]), .B(
        b11_OFWNT9L_8tZ[134]), .C(b4_nUAi[726]), .D(b4_nUAi[727]), .Y(
        b3_P_F_6_bm_230));
    
endmodule


module b8_1LbcQDr1_x_273_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [103:103] mdiclink_reg;
input  [273:273] b11_OFWNT9L_8tZ;
input  [311:309] b4_nUAi;
output [103:103] b6_2ZTGIf;

    wire b3_P_F_6_bm_2, b3_P_F_6_am_2, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_2), .B(
        b4_nUAi[311]), .C(b3_P_F_6_am_2), .Y(b6_2ZTGIf[103]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[103]), .B(
        b11_OFWNT9L_8tZ[273]), .C(b4_nUAi[310]), .D(b4_nUAi[309]), .Y(
        b3_P_F_6_am_2));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[103]), .B(
        b11_OFWNT9L_8tZ[273]), .C(b4_nUAi[309]), .D(b4_nUAi[310]), .Y(
        b3_P_F_6_bm_2));
    
endmodule


module b8_1LbcQDr1_x_320_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [56:56] mdiclink_reg;
input  [320:320] b11_OFWNT9L_8tZ;
input  [170:168] b4_nUAi;
output [56:56] b6_2ZTGIf;

    wire b3_P_F_6_bm_185, b3_P_F_6_am_185, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_185), .B(
        b4_nUAi[170]), .C(b3_P_F_6_am_185), .Y(b6_2ZTGIf[56]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[56]), .B(
        b11_OFWNT9L_8tZ[320]), .C(b4_nUAi[169]), .D(b4_nUAi[168]), .Y(
        b3_P_F_6_am_185));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[56]), .B(
        b11_OFWNT9L_8tZ[320]), .C(b4_nUAi[168]), .D(b4_nUAi[169]), .Y(
        b3_P_F_6_bm_185));
    
endmodule


module b8_1LbcQDr1_x_121_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [255:255] mdiclink_reg;
input  [121:121] b11_OFWNT9L_8tZ;
input  [766:765] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[255]), .B(
        b11_OFWNT9L_8tZ[121]), .C(b4_nUAi[766]), .D(b4_nUAi[765]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[255]), .B(
        b11_OFWNT9L_8tZ[121]), .C(b4_nUAi[766]), .D(b4_nUAi[765]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_142_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [234:234] mdiclink_reg;
input  [142:142] b11_OFWNT9L_8tZ;
input  [704:702] b4_nUAi;
output [234:234] b6_2ZTGIf;

    wire b3_P_F_6_bm_213, b3_P_F_6_am_213, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_213), .B(
        b4_nUAi[704]), .C(b3_P_F_6_am_213), .Y(b6_2ZTGIf[234]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[234]), .B(
        b11_OFWNT9L_8tZ[142]), .C(b4_nUAi[703]), .D(b4_nUAi[702]), .Y(
        b3_P_F_6_am_213));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[234]), .B(
        b11_OFWNT9L_8tZ[142]), .C(b4_nUAi[702]), .D(b4_nUAi[703]), .Y(
        b3_P_F_6_bm_213));
    
endmodule


module b8_1LbcQDr1_x_186_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [190:190] mdiclink_reg;
input  [186:186] b11_OFWNT9L_8tZ;
input  [571:570] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[190]), .B(
        b11_OFWNT9L_8tZ[186]), .C(b4_nUAi[571]), .D(b4_nUAi[570]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[190]), .B(
        b11_OFWNT9L_8tZ[186]), .C(b4_nUAi[571]), .D(b4_nUAi[570]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_292_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [84:84] mdiclink_reg;
input  [292:292] b11_OFWNT9L_8tZ;
input  [254:252] b4_nUAi;
output [84:84] b6_2ZTGIf;

    wire b3_P_F_6_bm_208, b3_P_F_6_am_208, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_208), .B(
        b4_nUAi[254]), .C(b3_P_F_6_am_208), .Y(b6_2ZTGIf[84]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[84]), .B(
        b11_OFWNT9L_8tZ[292]), .C(b4_nUAi[253]), .D(b4_nUAi[252]), .Y(
        b3_P_F_6_am_208));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[84]), .B(
        b11_OFWNT9L_8tZ[292]), .C(b4_nUAi[252]), .D(b4_nUAi[253]), .Y(
        b3_P_F_6_bm_208));
    
endmodule


module b8_1LbcQDr1_x_224_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [152:152] mdiclink_reg;
input  [224:224] b11_OFWNT9L_8tZ;
input  [458:456] b4_nUAi;
output [152:152] b6_2ZTGIf;

    wire b3_P_F_6_bm_31, b3_P_F_6_am_31, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_31), .B(
        b4_nUAi[458]), .C(b3_P_F_6_am_31), .Y(b6_2ZTGIf[152]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[152]), .B(
        b11_OFWNT9L_8tZ[224]), .C(b4_nUAi[457]), .D(b4_nUAi[456]), .Y(
        b3_P_F_6_am_31));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[152]), .B(
        b11_OFWNT9L_8tZ[224]), .C(b4_nUAi[456]), .D(b4_nUAi[457]), .Y(
        b3_P_F_6_bm_31));
    
endmodule


module b8_1LbcQDr1_x_195_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [181:181] mdiclink_reg;
input  [195:195] b11_OFWNT9L_8tZ;
input  [544:543] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[181]), .B(
        b11_OFWNT9L_8tZ[195]), .C(b4_nUAi[544]), .D(b4_nUAi[543]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[181]), .B(
        b11_OFWNT9L_8tZ[195]), .C(b4_nUAi[544]), .D(b4_nUAi[543]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_53_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [323:323] mdiclink_reg;
input  [53:53] b11_OFWNT9L_8tZ;
input  [971:969] b4_nUAi;
output [323:323] b6_2ZTGIf;

    wire b3_P_F_6_bm_125, b3_P_F_6_am_125, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_125), .B(
        b4_nUAi[971]), .C(b3_P_F_6_am_125), .Y(b6_2ZTGIf[323]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[323]), .B(
        b11_OFWNT9L_8tZ[53]), .C(b4_nUAi[970]), .D(b4_nUAi[969]), .Y(
        b3_P_F_6_am_125));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[323]), .B(
        b11_OFWNT9L_8tZ[53]), .C(b4_nUAi[969]), .D(b4_nUAi[970]), .Y(
        b3_P_F_6_bm_125));
    
endmodule


module b8_1LbcQDr1_x_15_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [361:361] mdiclink_reg;
input  [15:15] b11_OFWNT9L_8tZ;
input  [1085:1083] b4_nUAi;
output [361:361] b6_2ZTGIf;

    wire b3_P_F_6_bm_140, b3_P_F_6_am_140, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_140), .B(
        b4_nUAi[1085]), .C(b3_P_F_6_am_140), .Y(b6_2ZTGIf[361]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[361]), .B(
        b11_OFWNT9L_8tZ[15]), .C(b4_nUAi[1084]), .D(b4_nUAi[1083]), .Y(
        b3_P_F_6_am_140));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[361]), .B(
        b11_OFWNT9L_8tZ[15]), .C(b4_nUAi[1083]), .D(b4_nUAi[1084]), .Y(
        b3_P_F_6_bm_140));
    
endmodule


module b8_1LbcQDr1_x_100_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [276:276] mdiclink_reg;
input  [100:100] b11_OFWNT9L_8tZ;
input  [830:828] b4_nUAi;
output [276:276] b6_2ZTGIf;

    wire b3_P_F_6_bm_94, b3_P_F_6_am_94, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_94), .B(
        b4_nUAi[830]), .C(b3_P_F_6_am_94), .Y(b6_2ZTGIf[276]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[276]), .B(
        b11_OFWNT9L_8tZ[100]), .C(b4_nUAi[829]), .D(b4_nUAi[828]), .Y(
        b3_P_F_6_am_94));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[276]), .B(
        b11_OFWNT9L_8tZ[100]), .C(b4_nUAi[828]), .D(b4_nUAi[829]), .Y(
        b3_P_F_6_bm_94));
    
endmodule


module b8_1LbcQDr1_x_40_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [336:336] mdiclink_reg;
input  [40:40] b11_OFWNT9L_8tZ;
input  [1010:1008] b4_nUAi;
output [336:336] b6_2ZTGIf;

    wire b3_P_F_6_bm_138, b3_P_F_6_am_138, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_138), .B(
        b4_nUAi[1010]), .C(b3_P_F_6_am_138), .Y(b6_2ZTGIf[336]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[336]), .B(
        b11_OFWNT9L_8tZ[40]), .C(b4_nUAi[1009]), .D(b4_nUAi[1008]), .Y(
        b3_P_F_6_am_138));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[336]), .B(
        b11_OFWNT9L_8tZ[40]), .C(b4_nUAi[1008]), .D(b4_nUAi[1009]), .Y(
        b3_P_F_6_bm_138));
    
endmodule


module b8_1LbcQDr1_x_287_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [89:89] mdiclink_reg;
input  [287:287] b11_OFWNT9L_8tZ;
input  [269:267] b4_nUAi;
output [89:89] b6_2ZTGIf;

    wire b3_P_F_6_bm_204, b3_P_F_6_am_204, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_204), .B(
        b4_nUAi[269]), .C(b3_P_F_6_am_204), .Y(b6_2ZTGIf[89]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[89]), .B(
        b11_OFWNT9L_8tZ[287]), .C(b4_nUAi[268]), .D(b4_nUAi[267]), .Y(
        b3_P_F_6_am_204));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[89]), .B(
        b11_OFWNT9L_8tZ[287]), .C(b4_nUAi[267]), .D(b4_nUAi[268]), .Y(
        b3_P_F_6_bm_204));
    
endmodule


module b8_1LbcQDr1_x_35_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [341:341] mdiclink_reg;
input  [35:35] b11_OFWNT9L_8tZ;
input  [1024:1023] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[341]), .B(
        b11_OFWNT9L_8tZ[35]), .C(b4_nUAi[1024]), .D(b4_nUAi[1023]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[341]), .B(
        b11_OFWNT9L_8tZ[35]), .C(b4_nUAi[1024]), .D(b4_nUAi[1023]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_185_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [191:191] mdiclink_reg;
input  [185:185] b11_OFWNT9L_8tZ;
input  [574:573] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[191]), .B(
        b11_OFWNT9L_8tZ[185]), .C(b4_nUAi[574]), .D(b4_nUAi[573]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[191]), .B(
        b11_OFWNT9L_8tZ[185]), .C(b4_nUAi[574]), .D(b4_nUAi[573]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_375_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [1:1] mdiclink_reg;
input  [375:375] b11_OFWNT9L_8tZ;
input  [5:3] b4_nUAi;
output [1:1] b6_2ZTGIf;

    wire b3_P_F_6_bm_161, b3_P_F_6_am_161, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_161), .B(
        b4_nUAi[5]), .C(b3_P_F_6_am_161), .Y(b6_2ZTGIf[1]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[1]), .B(
        b11_OFWNT9L_8tZ[375]), .C(b4_nUAi[4]), .D(b4_nUAi[3]), .Y(
        b3_P_F_6_am_161));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[1]), .B(
        b11_OFWNT9L_8tZ[375]), .C(b4_nUAi[3]), .D(b4_nUAi[4]), .Y(
        b3_P_F_6_bm_161));
    
endmodule


module b8_1LbcQDr1_x_113_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [263:263] mdiclink_reg;
input  [113:113] b11_OFWNT9L_8tZ;
input  [791:789] b4_nUAi;
output [263:263] b6_2ZTGIf;

    wire b3_P_F_6_bm_82, b3_P_F_6_am_82, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_82), .B(
        b4_nUAi[791]), .C(b3_P_F_6_am_82), .Y(b6_2ZTGIf[263]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[263]), .B(
        b11_OFWNT9L_8tZ[113]), .C(b4_nUAi[790]), .D(b4_nUAi[789]), .Y(
        b3_P_F_6_am_82));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[263]), .B(
        b11_OFWNT9L_8tZ[113]), .C(b4_nUAi[789]), .D(b4_nUAi[790]), .Y(
        b3_P_F_6_bm_82));
    
endmodule


module b8_1LbcQDr1_x_221_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [155:155] mdiclink_reg;
input  [221:221] b11_OFWNT9L_8tZ;
input  [466:465] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[155]), .B(
        b11_OFWNT9L_8tZ[221]), .C(b4_nUAi[466]), .D(b4_nUAi[465]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[155]), .B(
        b11_OFWNT9L_8tZ[221]), .C(b4_nUAi[466]), .D(b4_nUAi[465]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_282_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [94:94] mdiclink_reg;
input  [282:282] b11_OFWNT9L_8tZ;
input  [283:282] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[94]), .B(
        b11_OFWNT9L_8tZ[282]), .C(b4_nUAi[283]), .D(b4_nUAi[282]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[94]), .B(
        b11_OFWNT9L_8tZ[282]), .C(b4_nUAi[283]), .D(b4_nUAi[282]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_151_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [225:225] mdiclink_reg;
input  [151:151] b11_OFWNT9L_8tZ;
input  [677:675] b4_nUAi;
output [225:225] b6_2ZTGIf;

    wire b3_P_F_6_bm_221, b3_P_F_6_am_221, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_221), .B(
        b4_nUAi[677]), .C(b3_P_F_6_am_221), .Y(b6_2ZTGIf[225]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[225]), .B(
        b11_OFWNT9L_8tZ[151]), .C(b4_nUAi[676]), .D(b4_nUAi[675]), .Y(
        b3_P_F_6_am_221));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[225]), .B(
        b11_OFWNT9L_8tZ[151]), .C(b4_nUAi[675]), .D(b4_nUAi[676]), .Y(
        b3_P_F_6_bm_221));
    
endmodule


module b8_1LbcQDr1_x_254_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [122:122] mdiclink_reg;
input  [254:254] b11_OFWNT9L_8tZ;
input  [368:366] b4_nUAi;
output [122:122] b6_2ZTGIf;

    wire b3_P_F_6_bm_9, b3_P_F_6_am_9, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_9), .B(
        b4_nUAi[368]), .C(b3_P_F_6_am_9), .Y(b6_2ZTGIf[122]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[122]), .B(
        b11_OFWNT9L_8tZ[254]), .C(b4_nUAi[367]), .D(b4_nUAi[366]), .Y(
        b3_P_F_6_am_9));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[122]), .B(
        b11_OFWNT9L_8tZ[254]), .C(b4_nUAi[366]), .D(b4_nUAi[367]), .Y(
        b3_P_F_6_bm_9));
    
endmodule


module b8_1LbcQDr1_x_39_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [337:337] mdiclink_reg;
input  [39:39] b11_OFWNT9L_8tZ;
input  [1013:1011] b4_nUAi;
output [337:337] b6_2ZTGIf;

    wire b3_P_F_6_bm_137, b3_P_F_6_am_137, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_137), .B(
        b4_nUAi[1013]), .C(b3_P_F_6_am_137), .Y(b6_2ZTGIf[337]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[337]), .B(
        b11_OFWNT9L_8tZ[39]), .C(b4_nUAi[1012]), .D(b4_nUAi[1011]), .Y(
        b3_P_F_6_am_137));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[337]), .B(
        b11_OFWNT9L_8tZ[39]), .C(b4_nUAi[1011]), .D(b4_nUAi[1012]), .Y(
        b3_P_F_6_bm_137));
    
endmodule


module b8_1LbcQDr1_x_367_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [9:9] mdiclink_reg;
input  [367:367] b11_OFWNT9L_8tZ;
input  [29:27] b4_nUAi;
output [9:9] b6_2ZTGIf;

    wire b3_P_F_6_bm_154, b3_P_F_6_am_154, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_154), .B(
        b4_nUAi[29]), .C(b3_P_F_6_am_154), .Y(b6_2ZTGIf[9]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[9]), .B(
        b11_OFWNT9L_8tZ[367]), .C(b4_nUAi[28]), .D(b4_nUAi[27]), .Y(
        b3_P_F_6_am_154));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[9]), .B(
        b11_OFWNT9L_8tZ[367]), .C(b4_nUAi[27]), .D(b4_nUAi[28]), .Y(
        b3_P_F_6_bm_154));
    
endmodule


module b8_1LbcQDr1_x_133_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [243:243] mdiclink_reg;
input  [133:133] b11_OFWNT9L_8tZ;
input  [731:729] b4_nUAi;
output [243:243] b6_2ZTGIf;

    wire b3_P_F_6_bm_229, b3_P_F_6_am_229, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_229), .B(
        b4_nUAi[731]), .C(b3_P_F_6_am_229), .Y(b6_2ZTGIf[243]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[243]), .B(
        b11_OFWNT9L_8tZ[133]), .C(b4_nUAi[730]), .D(b4_nUAi[729]), .Y(
        b3_P_F_6_am_229));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[243]), .B(
        b11_OFWNT9L_8tZ[133]), .C(b4_nUAi[729]), .D(b4_nUAi[730]), .Y(
        b3_P_F_6_bm_229));
    
endmodule


module b8_1LbcQDr1_x_162_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [214:214] mdiclink_reg;
input  [162:162] b11_OFWNT9L_8tZ;
input  [644:642] b4_nUAi;
output [214:214] b6_2ZTGIf;

    wire b3_P_F_6_bm_73, b3_P_F_6_am_73, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_73), .B(
        b4_nUAi[644]), .C(b3_P_F_6_am_73), .Y(b6_2ZTGIf[214]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[214]), .B(
        b11_OFWNT9L_8tZ[162]), .C(b4_nUAi[643]), .D(b4_nUAi[642]), .Y(
        b3_P_F_6_am_73));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[214]), .B(
        b11_OFWNT9L_8tZ[162]), .C(b4_nUAi[642]), .D(b4_nUAi[643]), .Y(
        b3_P_F_6_bm_73));
    
endmodule


module b8_1LbcQDr1_x_217_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [159:159] mdiclink_reg;
input  [217:217] b11_OFWNT9L_8tZ;
input  [478:477] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[159]), .B(
        b11_OFWNT9L_8tZ[217]), .C(b4_nUAi[478]), .D(b4_nUAi[477]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[159]), .B(
        b11_OFWNT9L_8tZ[217]), .C(b4_nUAi[478]), .D(b4_nUAi[477]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_172_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [204:204] mdiclink_reg;
input  [172:172] b11_OFWNT9L_8tZ;
input  [613:612] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[204]), .B(
        b11_OFWNT9L_8tZ[172]), .C(b4_nUAi[613]), .D(b4_nUAi[612]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[204]), .B(
        b11_OFWNT9L_8tZ[172]), .C(b4_nUAi[613]), .D(b4_nUAi[612]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_348_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [28:28] mdiclink_reg;
input  [348:348] b11_OFWNT9L_8tZ;
input  [85:84] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[28]), .B(
        b11_OFWNT9L_8tZ[348]), .C(b4_nUAi[85]), .D(b4_nUAi[84]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[28]), .B(
        b11_OFWNT9L_8tZ[348]), .C(b4_nUAi[85]), .D(b4_nUAi[84]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_144_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [232:232] mdiclink_reg;
input  [144:144] b11_OFWNT9L_8tZ;
input  [698:696] b4_nUAi;
output [232:232] b6_2ZTGIf;

    wire b3_P_F_6_bm_215, b3_P_F_6_am_215, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_215), .B(
        b4_nUAi[698]), .C(b3_P_F_6_am_215), .Y(b6_2ZTGIf[232]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[232]), .B(
        b11_OFWNT9L_8tZ[144]), .C(b4_nUAi[697]), .D(b4_nUAi[696]), .Y(
        b3_P_F_6_am_215));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[232]), .B(
        b11_OFWNT9L_8tZ[144]), .C(b4_nUAi[696]), .D(b4_nUAi[697]), .Y(
        b3_P_F_6_bm_215));
    
endmodule


module b8_1LbcQDr1_x_218_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [158:158] mdiclink_reg;
input  [218:218] b11_OFWNT9L_8tZ;
input  [475:474] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[158]), .B(
        b11_OFWNT9L_8tZ[218]), .C(b4_nUAi[475]), .D(b4_nUAi[474]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[158]), .B(
        b11_OFWNT9L_8tZ[218]), .C(b4_nUAi[475]), .D(b4_nUAi[474]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_308_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [68:68] mdiclink_reg;
input  [308:308] b11_OFWNT9L_8tZ;
input  [206:204] b4_nUAi;
output [68:68] b6_2ZTGIf;

    wire b3_P_F_6_bm_198, b3_P_F_6_am_198, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_198), .B(
        b4_nUAi[206]), .C(b3_P_F_6_am_198), .Y(b6_2ZTGIf[68]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[68]), .B(
        b11_OFWNT9L_8tZ[308]), .C(b4_nUAi[205]), .D(b4_nUAi[204]), .Y(
        b3_P_F_6_am_198));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[68]), .B(
        b11_OFWNT9L_8tZ[308]), .C(b4_nUAi[204]), .D(b4_nUAi[205]), .Y(
        b3_P_F_6_bm_198));
    
endmodule


module b8_1LbcQDr1_x_279_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [97:97] mdiclink_reg;
input  [279:279] b11_OFWNT9L_8tZ;
input  [293:291] b4_nUAi;
output [97:97] b6_2ZTGIf;

    wire b3_P_F_6_bm_7, b3_P_F_6_am_7, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_7), .B(
        b4_nUAi[293]), .C(b3_P_F_6_am_7), .Y(b6_2ZTGIf[97]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[97]), .B(
        b11_OFWNT9L_8tZ[279]), .C(b4_nUAi[292]), .D(b4_nUAi[291]), .Y(
        b3_P_F_6_am_7));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[97]), .B(
        b11_OFWNT9L_8tZ[279]), .C(b4_nUAi[291]), .D(b4_nUAi[292]), .Y(
        b3_P_F_6_bm_7));
    
endmodule


module b8_1LbcQDr1_x_60_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [316:316] mdiclink_reg;
input  [60:60] b11_OFWNT9L_8tZ;
input  [949:948] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[316]), .B(
        b11_OFWNT9L_8tZ[60]), .C(b4_nUAi[949]), .D(b4_nUAi[948]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[316]), .B(
        b11_OFWNT9L_8tZ[60]), .C(b4_nUAi[949]), .D(b4_nUAi[948]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_303_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [73:73] mdiclink_reg;
input  [303:303] b11_OFWNT9L_8tZ;
input  [221:219] b4_nUAi;
output [73:73] b6_2ZTGIf;

    wire b3_P_F_6_bm_194, b3_P_F_6_am_194, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_194), .B(
        b4_nUAi[221]), .C(b3_P_F_6_am_194), .Y(b6_2ZTGIf[73]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[73]), .B(
        b11_OFWNT9L_8tZ[303]), .C(b4_nUAi[220]), .D(b4_nUAi[219]), .Y(
        b3_P_F_6_am_194));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[73]), .B(
        b11_OFWNT9L_8tZ[303]), .C(b4_nUAi[219]), .D(b4_nUAi[220]), .Y(
        b3_P_F_6_bm_194));
    
endmodule


module b8_1LbcQDr1_x_363_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [13:13] mdiclink_reg;
input  [363:363] b11_OFWNT9L_8tZ;
input  [40:39] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[13]), .B(
        b11_OFWNT9L_8tZ[363]), .C(b4_nUAi[40]), .D(b4_nUAi[39]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[13]), .B(
        b11_OFWNT9L_8tZ[363]), .C(b4_nUAi[40]), .D(b4_nUAi[39]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_108_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [268:268] mdiclink_reg;
input  [108:108] b11_OFWNT9L_8tZ;
input  [805:804] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[268]), .B(
        b11_OFWNT9L_8tZ[108]), .C(b4_nUAi[805]), .D(b4_nUAi[804]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[268]), .B(
        b11_OFWNT9L_8tZ[108]), .C(b4_nUAi[805]), .D(b4_nUAi[804]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_333_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [43:43] mdiclink_reg;
input  [333:333] b11_OFWNT9L_8tZ;
input  [130:129] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[43]), .B(
        b11_OFWNT9L_8tZ[333]), .C(b4_nUAi[130]), .D(b4_nUAi[129]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[43]), .B(
        b11_OFWNT9L_8tZ[333]), .C(b4_nUAi[130]), .D(b4_nUAi[129]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_219_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [157:157] mdiclink_reg;
input  [219:219] b11_OFWNT9L_8tZ;
input  [472:471] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[157]), .B(
        b11_OFWNT9L_8tZ[219]), .C(b4_nUAi[472]), .D(b4_nUAi[471]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[157]), .B(
        b11_OFWNT9L_8tZ[219]), .C(b4_nUAi[472]), .D(b4_nUAi[471]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_70_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [306:306] mdiclink_reg;
input  [70:70] b11_OFWNT9L_8tZ;
input  [920:918] b4_nUAi;
output [306:306] b6_2ZTGIf;

    wire b3_P_F_6_bm_116, b3_P_F_6_am_116, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_116), .B(
        b4_nUAi[920]), .C(b3_P_F_6_am_116), .Y(b6_2ZTGIf[306]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[306]), .B(
        b11_OFWNT9L_8tZ[70]), .C(b4_nUAi[919]), .D(b4_nUAi[918]), .Y(
        b3_P_F_6_am_116));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[306]), .B(
        b11_OFWNT9L_8tZ[70]), .C(b4_nUAi[918]), .D(b4_nUAi[919]), .Y(
        b3_P_F_6_bm_116));
    
endmodule


module b8_1LbcQDr1_x_251_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [125:125] mdiclink_reg;
input  [251:251] b11_OFWNT9L_8tZ;
input  [376:375] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[125]), .B(
        b11_OFWNT9L_8tZ[251]), .C(b4_nUAi[376]), .D(b4_nUAi[375]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[125]), .B(
        b11_OFWNT9L_8tZ[251]), .C(b4_nUAi[376]), .D(b4_nUAi[375]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_323_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [53:53] mdiclink_reg;
input  [323:323] b11_OFWNT9L_8tZ;
input  [160:159] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[53]), .B(
        b11_OFWNT9L_8tZ[323]), .C(b4_nUAi[160]), .D(b4_nUAi[159]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[53]), .B(
        b11_OFWNT9L_8tZ[323]), .C(b4_nUAi[160]), .D(b4_nUAi[159]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_95_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [281:281] mdiclink_reg;
input  [95:95] b11_OFWNT9L_8tZ;
input  [845:843] b4_nUAi;
output [281:281] b6_2ZTGIf;

    wire b3_P_F_6_bm_90, b3_P_F_6_am_90, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_90), .B(
        b4_nUAi[845]), .C(b3_P_F_6_am_90), .Y(b6_2ZTGIf[281]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[281]), .B(
        b11_OFWNT9L_8tZ[95]), .C(b4_nUAi[844]), .D(b4_nUAi[843]), .Y(
        b3_P_F_6_am_90));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[281]), .B(
        b11_OFWNT9L_8tZ[95]), .C(b4_nUAi[843]), .D(b4_nUAi[844]), .Y(
        b3_P_F_6_bm_90));
    
endmodule


module b8_1LbcQDr1_x_347_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [29:29] mdiclink_reg;
input  [347:347] b11_OFWNT9L_8tZ;
input  [88:87] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[29]), .B(
        b11_OFWNT9L_8tZ[347]), .C(b4_nUAi[88]), .D(b4_nUAi[87]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[29]), .B(
        b11_OFWNT9L_8tZ[347]), .C(b4_nUAi[88]), .D(b4_nUAi[87]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_226_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [150:150] mdiclink_reg;
input  [226:226] b11_OFWNT9L_8tZ;
input  [452:450] b4_nUAi;
output [150:150] b6_2ZTGIf;

    wire b3_P_F_6_bm_33, b3_P_F_6_am_33, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_33), .B(
        b4_nUAi[452]), .C(b3_P_F_6_am_33), .Y(b6_2ZTGIf[150]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[150]), .B(
        b11_OFWNT9L_8tZ[226]), .C(b4_nUAi[451]), .D(b4_nUAi[450]), .Y(
        b3_P_F_6_am_33));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[150]), .B(
        b11_OFWNT9L_8tZ[226]), .C(b4_nUAi[450]), .D(b4_nUAi[451]), .Y(
        b3_P_F_6_bm_33));
    
endmodule


module b8_1LbcQDr1_x_128_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [248:248] mdiclink_reg;
input  [128:128] b11_OFWNT9L_8tZ;
input  [746:744] b4_nUAi;
output [248:248] b6_2ZTGIf;

    wire b3_P_F_6_bm_225, b3_P_F_6_am_225, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_225), .B(
        b4_nUAi[746]), .C(b3_P_F_6_am_225), .Y(b6_2ZTGIf[248]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[248]), .B(
        b11_OFWNT9L_8tZ[128]), .C(b4_nUAi[745]), .D(b4_nUAi[744]), .Y(
        b3_P_F_6_am_225));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[248]), .B(
        b11_OFWNT9L_8tZ[128]), .C(b4_nUAi[744]), .D(b4_nUAi[745]), .Y(
        b3_P_F_6_bm_225));
    
endmodule


module b8_1LbcQDr1_x_307_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [69:69] mdiclink_reg;
input  [307:307] b11_OFWNT9L_8tZ;
input  [208:207] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[69]), .B(
        b11_OFWNT9L_8tZ[307]), .C(b4_nUAi[208]), .D(b4_nUAi[207]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[69]), .B(
        b11_OFWNT9L_8tZ[307]), .C(b4_nUAi[208]), .D(b4_nUAi[207]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_330_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [46:46] mdiclink_reg;
input  [330:330] b11_OFWNT9L_8tZ;
input  [139:138] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[46]), .B(
        b11_OFWNT9L_8tZ[330]), .C(b4_nUAi[139]), .D(b4_nUAi[138]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[46]), .B(
        b11_OFWNT9L_8tZ[330]), .C(b4_nUAi[139]), .D(b4_nUAi[138]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_12_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [364:364] mdiclink_reg;
input  [12:12] b11_OFWNT9L_8tZ;
input  [1093:1092] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[364]), .B(
        b11_OFWNT9L_8tZ[12]), .C(b4_nUAi[1093]), .D(b4_nUAi[1092]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[364]), .B(
        b11_OFWNT9L_8tZ[12]), .C(b4_nUAi[1093]), .D(b4_nUAi[1092]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_193_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [183:183] mdiclink_reg;
input  [193:193] b11_OFWNT9L_8tZ;
input  [551:549] b4_nUAi;
output [183:183] b6_2ZTGIf;

    wire b3_P_F_6_bm_52, b3_P_F_6_am_52, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_52), .B(
        b4_nUAi[551]), .C(b3_P_F_6_am_52), .Y(b6_2ZTGIf[183]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[183]), .B(
        b11_OFWNT9L_8tZ[193]), .C(b4_nUAi[550]), .D(b4_nUAi[549]), .Y(
        b3_P_F_6_am_52));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[183]), .B(
        b11_OFWNT9L_8tZ[193]), .C(b4_nUAi[549]), .D(b4_nUAi[550]), .Y(
        b3_P_F_6_bm_52));
    
endmodule


module b8_1LbcQDr1_x_45_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [331:331] mdiclink_reg;
input  [45:45] b11_OFWNT9L_8tZ;
input  [994:993] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[331]), .B(
        b11_OFWNT9L_8tZ[45]), .C(b4_nUAi[994]), .D(b4_nUAi[993]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[331]), .B(
        b11_OFWNT9L_8tZ[45]), .C(b4_nUAi[994]), .D(b4_nUAi[993]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_21_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [355:355] mdiclink_reg;
input  [21:21] b11_OFWNT9L_8tZ;
input  [1067:1065] b4_nUAi;
output [355:355] b6_2ZTGIf;

    wire b3_P_F_6_bm_145, b3_P_F_6_am_145, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_145), .B(
        b4_nUAi[1067]), .C(b3_P_F_6_am_145), .Y(b6_2ZTGIf[355]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[355]), .B(
        b11_OFWNT9L_8tZ[21]), .C(b4_nUAi[1066]), .D(b4_nUAi[1065]), .Y(
        b3_P_F_6_am_145));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[355]), .B(
        b11_OFWNT9L_8tZ[21]), .C(b4_nUAi[1065]), .D(b4_nUAi[1066]), .Y(
        b3_P_F_6_bm_145));
    
endmodule


module b8_1LbcQDr1_x_3_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [373:373] mdiclink_reg;
input  [3:3] b11_OFWNT9L_8tZ;
input  [1121:1119] b4_nUAi;
output [373:373] b6_2ZTGIf;

    wire b3_P_F_6_bm_150, b3_P_F_6_am_150, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_150), .B(
        b4_nUAi[1121]), .C(b3_P_F_6_am_150), .Y(b6_2ZTGIf[373]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[373]), .B(
        b11_OFWNT9L_8tZ[3]), .C(b4_nUAi[1120]), .D(b4_nUAi[1119]), .Y(
        b3_P_F_6_am_150));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[373]), .B(
        b11_OFWNT9L_8tZ[3]), .C(b4_nUAi[1119]), .D(b4_nUAi[1120]), .Y(
        b3_P_F_6_bm_150));
    
endmodule


module b8_1LbcQDr1_x_116_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [260:260] mdiclink_reg;
input  [116:116] b11_OFWNT9L_8tZ;
input  [782:780] b4_nUAi;
output [260:260] b6_2ZTGIf;

    wire b3_P_F_6_bm_84, b3_P_F_6_am_84, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_84), .B(
        b4_nUAi[782]), .C(b3_P_F_6_am_84), .Y(b6_2ZTGIf[260]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[260]), .B(
        b11_OFWNT9L_8tZ[116]), .C(b4_nUAi[781]), .D(b4_nUAi[780]), .Y(
        b3_P_F_6_am_84));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[260]), .B(
        b11_OFWNT9L_8tZ[116]), .C(b4_nUAi[780]), .D(b4_nUAi[781]), .Y(
        b3_P_F_6_bm_84));
    
endmodule


module b8_1LbcQDr1_x_247_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [129:129] mdiclink_reg;
input  [247:247] b11_OFWNT9L_8tZ;
input  [389:387] b4_nUAi;
output [129:129] b6_2ZTGIf;

    wire b3_P_F_6_bm_27, b3_P_F_6_am_27, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_27), .B(
        b4_nUAi[389]), .C(b3_P_F_6_am_27), .Y(b6_2ZTGIf[129]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[129]), .B(
        b11_OFWNT9L_8tZ[247]), .C(b4_nUAi[388]), .D(b4_nUAi[387]), .Y(
        b3_P_F_6_am_27));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[129]), .B(
        b11_OFWNT9L_8tZ[247]), .C(b4_nUAi[387]), .D(b4_nUAi[388]), .Y(
        b3_P_F_6_bm_27));
    
endmodule


module b8_1LbcQDr1_x_59_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [317:317] mdiclink_reg;
input  [59:59] b11_OFWNT9L_8tZ;
input  [952:951] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[317]), .B(
        b11_OFWNT9L_8tZ[59]), .C(b4_nUAi[952]), .D(b4_nUAi[951]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[317]), .B(
        b11_OFWNT9L_8tZ[59]), .C(b4_nUAi[952]), .D(b4_nUAi[951]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_291_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [85:85] mdiclink_reg;
input  [291:291] b11_OFWNT9L_8tZ;
input  [256:255] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[85]), .B(
        b11_OFWNT9L_8tZ[291]), .C(b4_nUAi[256]), .D(b4_nUAi[255]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[85]), .B(
        b11_OFWNT9L_8tZ[291]), .C(b4_nUAi[256]), .D(b4_nUAi[255]), .Y(
        N_25));
    
endmodule


module b11_PSyil9s1fkT_x(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b11_uUT0JC4gFrY,
       BW_clk_c,
       b7_PSyi3wy
    );
input  [376:0] mdiclink_reg;
input  [376:0] b11_OFWNT9L_8tZ;
input  [1129:0] b4_nUAi;
output [1:1] b11_uUT0JC4gFrY;
input  BW_clk_c;
input  b7_PSyi3wy;

    wire \b6_2ZTGIf[0] , \b6_2ZTGIf[1] , \b6_2ZTGIf[2] , 
        \b6_2ZTGIf[3] , \b6_2ZTGIf[4] , N_27, N_25, \b6_2ZTGIf[6] , 
        \b6_2ZTGIf[7] , \b6_2ZTGIf[8] , \b6_2ZTGIf[9] , 
        \b6_2ZTGIf[10] , N_27_0, N_25_0, N_27_1, N_25_1, N_27_2, 
        N_25_2, N_27_3, N_25_3, N_27_4, N_25_4, \b6_2ZTGIf[16] , 
        \b6_2ZTGIf[17] , \b6_2ZTGIf[18] , \b6_2ZTGIf[19] , 
        \b6_2ZTGIf[20] , N_27_5, N_25_5, \b6_2ZTGIf[22] , 
        \b6_2ZTGIf[23] , \b6_2ZTGIf[24] , \b6_2ZTGIf[25] , 
        \b6_2ZTGIf[26] , N_27_6, N_25_6, N_27_7, N_25_7, N_27_8, 
        N_25_8, N_27_9, N_25_9, N_27_10, N_25_10, \b6_2ZTGIf[32] , 
        \b6_2ZTGIf[33] , \b6_2ZTGIf[34] , \b6_2ZTGIf[35] , 
        \b6_2ZTGIf[36] , N_27_11, N_25_11, \b6_2ZTGIf[38] , 
        \b6_2ZTGIf[39] , \b6_2ZTGIf[40] , \b6_2ZTGIf[41] , 
        \b6_2ZTGIf[42] , N_27_12, N_25_12, N_27_13, N_25_13, N_27_14, 
        N_25_14, N_27_15, N_25_15, N_27_16, N_25_16, \b6_2ZTGIf[48] , 
        \b6_2ZTGIf[49] , \b6_2ZTGIf[50] , \b6_2ZTGIf[51] , 
        \b6_2ZTGIf[52] , N_27_17, N_25_17, \b6_2ZTGIf[54] , 
        \b6_2ZTGIf[55] , \b6_2ZTGIf[56] , \b6_2ZTGIf[57] , 
        \b6_2ZTGIf[58] , N_27_18, N_25_18, N_27_19, N_25_19, N_27_20, 
        N_25_20, N_27_21, N_25_21, N_27_22, N_25_22, \b6_2ZTGIf[64] , 
        \b6_2ZTGIf[65] , \b6_2ZTGIf[66] , \b6_2ZTGIf[67] , 
        \b6_2ZTGIf[68] , N_27_23, N_25_23, \b6_2ZTGIf[70] , 
        \b6_2ZTGIf[71] , \b6_2ZTGIf[72] , \b6_2ZTGIf[73] , 
        \b6_2ZTGIf[74] , N_27_24, N_25_24, N_27_25, N_25_25, N_27_26, 
        N_25_26, N_27_27, N_25_27, N_27_28, N_25_28, \b6_2ZTGIf[80] , 
        \b6_2ZTGIf[81] , \b6_2ZTGIf[82] , \b6_2ZTGIf[83] , 
        \b6_2ZTGIf[84] , N_27_29, N_25_29, \b6_2ZTGIf[86] , 
        \b6_2ZTGIf[87] , \b6_2ZTGIf[88] , \b6_2ZTGIf[89] , 
        \b6_2ZTGIf[90] , N_27_30, N_25_30, N_27_31, N_25_31, N_27_32, 
        N_25_32, N_27_33, N_25_33, N_27_34, N_25_34, \b6_2ZTGIf[96] , 
        \b6_2ZTGIf[97] , \b6_2ZTGIf[98] , \b6_2ZTGIf[99] , 
        \b6_2ZTGIf[100] , N_27_35, N_25_35, \b6_2ZTGIf[102] , 
        \b6_2ZTGIf[103] , \b6_2ZTGIf[104] , \b6_2ZTGIf[105] , 
        \b6_2ZTGIf[106] , N_27_36, N_25_36, N_27_37, N_25_37, N_27_38, 
        N_25_38, N_27_39, N_25_39, N_27_40, N_25_40, \b6_2ZTGIf[112] , 
        \b6_2ZTGIf[113] , \b6_2ZTGIf[114] , \b6_2ZTGIf[115] , 
        \b6_2ZTGIf[116] , N_27_41, N_25_41, \b6_2ZTGIf[118] , 
        \b6_2ZTGIf[119] , \b6_2ZTGIf[120] , \b6_2ZTGIf[121] , 
        \b6_2ZTGIf[122] , N_27_42, N_25_42, N_27_43, N_25_43, N_27_44, 
        N_25_44, N_27_45, N_25_45, N_27_46, N_25_46, \b6_2ZTGIf[128] , 
        \b6_2ZTGIf[129] , \b6_2ZTGIf[130] , \b6_2ZTGIf[131] , 
        \b6_2ZTGIf[132] , N_27_47, N_25_47, \b6_2ZTGIf[134] , 
        \b6_2ZTGIf[135] , \b6_2ZTGIf[136] , \b6_2ZTGIf[137] , 
        \b6_2ZTGIf[138] , N_27_48, N_25_48, N_27_49, N_25_49, N_27_50, 
        N_25_50, N_27_51, N_25_51, N_27_52, N_25_52, \b6_2ZTGIf[144] , 
        \b6_2ZTGIf[145] , \b6_2ZTGIf[146] , \b6_2ZTGIf[147] , 
        \b6_2ZTGIf[148] , N_27_53, N_25_53, \b6_2ZTGIf[150] , 
        \b6_2ZTGIf[151] , \b6_2ZTGIf[152] , \b6_2ZTGIf[153] , 
        \b6_2ZTGIf[154] , N_27_54, N_25_54, N_27_55, N_25_55, N_27_56, 
        N_25_56, N_27_57, N_25_57, N_27_58, N_25_58, \b6_2ZTGIf[160] , 
        \b6_2ZTGIf[161] , \b6_2ZTGIf[162] , \b6_2ZTGIf[163] , 
        \b6_2ZTGIf[164] , N_27_59, N_25_59, \b6_2ZTGIf[166] , 
        \b6_2ZTGIf[167] , \b6_2ZTGIf[168] , \b6_2ZTGIf[169] , 
        \b6_2ZTGIf[170] , N_27_60, N_25_60, N_27_61, N_25_61, N_27_62, 
        N_25_62, N_27_63, N_25_63, N_27_64, N_25_64, \b6_2ZTGIf[176] , 
        \b6_2ZTGIf[177] , \b6_2ZTGIf[178] , \b6_2ZTGIf[179] , 
        \b6_2ZTGIf[180] , N_27_65, N_25_65, \b6_2ZTGIf[182] , 
        \b6_2ZTGIf[183] , \b6_2ZTGIf[184] , \b6_2ZTGIf[185] , 
        \b6_2ZTGIf[186] , N_27_66, N_25_66, N_27_67, N_25_67, N_27_68, 
        N_25_68, N_27_69, N_25_69, N_27_70, N_25_70, \b6_2ZTGIf[192] , 
        \b6_2ZTGIf[193] , \b6_2ZTGIf[194] , \b6_2ZTGIf[195] , 
        \b6_2ZTGIf[196] , N_27_71, N_25_71, \b6_2ZTGIf[198] , 
        \b6_2ZTGIf[199] , \b6_2ZTGIf[200] , \b6_2ZTGIf[201] , 
        \b6_2ZTGIf[202] , N_27_72, N_25_72, N_27_73, N_25_73, N_27_74, 
        N_25_74, N_27_75, N_25_75, N_27_76, N_25_76, \b6_2ZTGIf[208] , 
        \b6_2ZTGIf[209] , \b6_2ZTGIf[210] , \b6_2ZTGIf[211] , 
        \b6_2ZTGIf[212] , N_27_77, N_25_77, \b6_2ZTGIf[214] , 
        \b6_2ZTGIf[215] , \b6_2ZTGIf[216] , \b6_2ZTGIf[217] , 
        \b6_2ZTGIf[218] , N_27_78, N_25_78, N_27_79, N_25_79, N_27_80, 
        N_25_80, N_27_81, N_25_81, N_27_82, N_25_82, \b6_2ZTGIf[224] , 
        \b6_2ZTGIf[225] , \b6_2ZTGIf[226] , \b6_2ZTGIf[227] , 
        \b6_2ZTGIf[228] , N_27_83, N_25_83, \b6_2ZTGIf[230] , 
        \b6_2ZTGIf[231] , \b6_2ZTGIf[232] , \b6_2ZTGIf[233] , 
        \b6_2ZTGIf[234] , N_27_84, N_25_84, N_27_85, N_25_85, N_27_86, 
        N_25_86, N_27_87, N_25_87, N_27_88, N_25_88, \b6_2ZTGIf[240] , 
        \b6_2ZTGIf[241] , \b6_2ZTGIf[242] , \b6_2ZTGIf[243] , 
        \b6_2ZTGIf[244] , N_27_89, N_25_89, \b6_2ZTGIf[246] , 
        \b6_2ZTGIf[247] , \b6_2ZTGIf[248] , \b6_2ZTGIf[249] , 
        \b6_2ZTGIf[250] , N_27_90, N_25_90, N_27_91, N_25_91, N_27_92, 
        N_25_92, N_27_93, N_25_93, N_27_94, N_25_94, \b6_2ZTGIf[256] , 
        \b6_2ZTGIf[257] , \b6_2ZTGIf[258] , \b6_2ZTGIf[259] , 
        \b6_2ZTGIf[260] , N_27_95, N_25_95, \b6_2ZTGIf[262] , 
        \b6_2ZTGIf[263] , \b6_2ZTGIf[264] , \b6_2ZTGIf[265] , 
        \b6_2ZTGIf[266] , N_27_96, N_25_96, N_27_97, N_25_97, N_27_98, 
        N_25_98, N_27_99, N_25_99, N_27_100, N_25_100, 
        \b6_2ZTGIf[272] , \b6_2ZTGIf[273] , \b6_2ZTGIf[274] , 
        \b6_2ZTGIf[275] , \b6_2ZTGIf[276] , N_27_101, N_25_101, 
        \b6_2ZTGIf[278] , \b6_2ZTGIf[279] , \b6_2ZTGIf[280] , 
        \b6_2ZTGIf[281] , \b6_2ZTGIf[282] , N_27_102, N_25_102, 
        N_27_103, N_25_103, N_27_104, N_25_104, N_27_105, N_25_105, 
        N_27_106, N_25_106, \b6_2ZTGIf[288] , \b6_2ZTGIf[289] , 
        \b6_2ZTGIf[290] , \b6_2ZTGIf[291] , \b6_2ZTGIf[292] , N_27_107, 
        N_25_107, \b6_2ZTGIf[294] , \b6_2ZTGIf[295] , \b6_2ZTGIf[296] , 
        \b6_2ZTGIf[297] , \b6_2ZTGIf[298] , N_27_108, N_25_108, 
        N_27_109, N_25_109, N_27_110, N_25_110, N_27_111, N_25_111, 
        N_27_112, N_25_112, \b6_2ZTGIf[304] , \b6_2ZTGIf[305] , 
        \b6_2ZTGIf[306] , \b6_2ZTGIf[307] , \b6_2ZTGIf[308] , N_27_113, 
        N_25_113, \b6_2ZTGIf[310] , \b6_2ZTGIf[311] , \b6_2ZTGIf[312] , 
        \b6_2ZTGIf[313] , \b6_2ZTGIf[314] , N_27_114, N_25_114, 
        N_27_115, N_25_115, N_27_116, N_25_116, N_27_117, N_25_117, 
        N_27_118, N_25_118, \b6_2ZTGIf[320] , \b6_2ZTGIf[321] , 
        \b6_2ZTGIf[322] , \b6_2ZTGIf[323] , \b6_2ZTGIf[324] , N_27_119, 
        N_25_119, \b6_2ZTGIf[326] , \b6_2ZTGIf[327] , \b6_2ZTGIf[328] , 
        \b6_2ZTGIf[329] , \b6_2ZTGIf[330] , N_27_120, N_25_120, 
        N_27_121, N_25_121, N_27_122, N_25_122, N_27_123, N_25_123, 
        N_27_124, N_25_124, \b6_2ZTGIf[336] , \b6_2ZTGIf[337] , 
        \b6_2ZTGIf[338] , \b6_2ZTGIf[339] , \b6_2ZTGIf[340] , N_27_125, 
        N_25_125, \b6_2ZTGIf[342] , \b6_2ZTGIf[343] , \b6_2ZTGIf[344] , 
        \b6_2ZTGIf[345] , \b6_2ZTGIf[346] , N_27_126, N_25_126, 
        N_27_127, N_25_127, N_27_128, N_25_128, N_27_129, N_25_129, 
        N_27_130, N_25_130, \b6_2ZTGIf[352] , \b6_2ZTGIf[353] , 
        \b6_2ZTGIf[354] , \b6_2ZTGIf[355] , \b6_2ZTGIf[356] , N_27_131, 
        N_25_131, \b6_2ZTGIf[358] , \b6_2ZTGIf[359] , \b6_2ZTGIf[360] , 
        \b6_2ZTGIf[361] , \b6_2ZTGIf[362] , N_27_132, N_25_132, 
        N_27_133, N_25_133, N_27_134, N_25_134, N_27_135, N_25_135, 
        N_27_136, N_25_136, N_27_137, N_25_137, \b6_2ZTGIf[369] , 
        N_27_138, N_25_138, \b6_2ZTGIf[371] , N_27_139, N_25_139, 
        \b6_2ZTGIf[373] , N_27_140, N_25_140, \b6_2ZTGIf[375] , 
        N_27_141, N_25_141, GND_net_1, VCC_net_1;
    
    b8_1LbcQDr1_x_85_0 b9_1LbcgKwVn (.mdiclink_reg({mdiclink_reg[291]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[85]}), .b4_nUAi({
        b4_nUAi[875], b4_nUAi[874], b4_nUAi[873]}), .b6_2ZTGIf({
        \b6_2ZTGIf[291] }));
    b8_1LbcQDr1_x_69_0 b9_1LbcgKeRe (.mdiclink_reg({mdiclink_reg[307]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[69]}), .b4_nUAi({
        b4_nUAi[923], b4_nUAi[922], b4_nUAi[921]}), .b6_2ZTGIf({
        \b6_2ZTGIf[307] }));
    b8_1LbcQDr1_x_16_0 b9_1LbcgKeAm (.mdiclink_reg({mdiclink_reg[360]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[16]}), .b4_nUAi({
        b4_nUAi[1082], b4_nUAi[1081], b4_nUAi[1080]}), .b6_2ZTGIf({
        \b6_2ZTGIf[360] }));
    b8_1LbcQDr1_x_248_0 b9_1LbcgKGIS (.mdiclink_reg({mdiclink_reg[128]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[248]}), .b4_nUAi({
        b4_nUAi[386], b4_nUAi[385], b4_nUAi[384]}), .b6_2ZTGIf({
        \b6_2ZTGIf[128] }));
    b8_1LbcQDr1_x_32_0 b9_1LbcgKeQl0 (.mdiclink_reg({mdiclink_reg[344]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[32]}), .b4_nUAi({
        b4_nUAi[1034], b4_nUAi[1033], b4_nUAi[1032]}), .b6_2ZTGIf({
        \b6_2ZTGIf[344] }));
    b8_1LbcQDr1_x_302_0 b8_1LbcgKxQ0 (.mdiclink_reg({mdiclink_reg[74]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[302]}), .b4_nUAi({
        b4_nUAi[224], b4_nUAi[223], b4_nUAi[222]}), .b6_2ZTGIf({
        \b6_2ZTGIf[74] }));
    b8_1LbcQDr1_x_136_0 b9_1LbcgKwQm0 (.mdiclink_reg({
        mdiclink_reg[240]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[136]}), 
        .b4_nUAi({b4_nUAi[722], b4_nUAi[721], b4_nUAi[720]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[240] }));
    b8_1LbcQDr1_x_225_0 b9_1LbcgKGUn (.mdiclink_reg({mdiclink_reg[151]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[225]}), .b4_nUAi({
        b4_nUAi[455], b4_nUAi[454], b4_nUAi[453]}), .b6_2ZTGIf({
        \b6_2ZTGIf[151] }));
    b8_1LbcQDr1_x_183_0 b9_1LbcgKGVV (.mdiclink_reg({mdiclink_reg[193]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[183]}), .b4_nUAi({
        b4_nUAi[581], b4_nUAi[580], b4_nUAi[579]}), .b6_2ZTGIf({
        \b6_2ZTGIf[193] }));
    b8_1LbcQDr1_x_249_0 b9_1LbcgKGIe (.mdiclink_reg({mdiclink_reg[127]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[249]}), .b4_nUAi({
        b4_nUAi[382], b4_nUAi[381]}), .N_27(N_27_46), .N_25(N_25_46));
    b8_1LbcQDr1_x_362_0 b8_1LbcgKGQ0 (.mdiclink_reg({mdiclink_reg[14]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[362]}), .b4_nUAi({
        b4_nUAi[43], b4_nUAi[42]}), .N_27(N_27_3), .N_25(N_25_3));
    b8_1LbcQDr1_x_164_0 b9_1LbcgKwSd (.mdiclink_reg({mdiclink_reg[212]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[164]}), .b4_nUAi({
        b4_nUAi[638], b4_nUAi[637], b4_nUAi[636]}), .b6_2ZTGIf({
        \b6_2ZTGIf[212] }));
    b8_1LbcQDr1_x_143_0 b9_1LbcgKwqV (.mdiclink_reg({mdiclink_reg[233]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[143]}), .b4_nUAi({
        b4_nUAi[701], b4_nUAi[700], b4_nUAi[699]}), .b6_2ZTGIf({
        \b6_2ZTGIf[233] }));
    b8_1LbcQDr1_x_36_0 b9_1LbcgKeQm0 (.mdiclink_reg({mdiclink_reg[340]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[36]}), .b4_nUAi({
        b4_nUAi[1022], b4_nUAi[1021], b4_nUAi[1020]}), .b6_2ZTGIf({
        \b6_2ZTGIf[340] }));
    b8_1LbcQDr1_x_24_0 b9_1LbcgKeUd (.mdiclink_reg({mdiclink_reg[352]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[24]}), .b4_nUAi({
        b4_nUAi[1058], b4_nUAi[1057], b4_nUAi[1056]}), .b6_2ZTGIf({
        \b6_2ZTGIf[352] }));
    b8_1LbcQDr1_x_174_0 b9_1LbcgKwRd (.mdiclink_reg({mdiclink_reg[202]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[174]}), .b4_nUAi({
        b4_nUAi[608], b4_nUAi[607], b4_nUAi[606]}), .b6_2ZTGIf({
        \b6_2ZTGIf[202] }));
    b8_1LbcQDr1_x_305_0 b8_1LbcgKxS (.mdiclink_reg({mdiclink_reg[71]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[305]}), .b4_nUAi({
        b4_nUAi[215], b4_nUAi[214], b4_nUAi[213]}), .b6_2ZTGIf({
        \b6_2ZTGIf[71] }));
    b8_1LbcQDr1_x_365_0 b8_1LbcgKGS (.mdiclink_reg({mdiclink_reg[11]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[365]}), .b4_nUAi({
        b4_nUAi[34], b4_nUAi[33]}), .N_27(N_27_0), .N_25(N_25_0));
    b8_1LbcQDr1_x_256_0 b9_1LbcgKGIm (.mdiclink_reg({mdiclink_reg[120]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[256]}), .b4_nUAi({
        b4_nUAi[362], b4_nUAi[361], b4_nUAi[360]}), .b6_2ZTGIf({
        \b6_2ZTGIf[120] }));
    b8_1LbcQDr1_x_101_0 b9_1LbcgKwJp (.mdiclink_reg({mdiclink_reg[275]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[101]}), .b4_nUAi({
        b4_nUAi[827], b4_nUAi[826], b4_nUAi[825]}), .b6_2ZTGIf({
        \b6_2ZTGIf[275] }));
    b8_1LbcQDr1_x_306_0 b8_1LbcgKxR (.mdiclink_reg({mdiclink_reg[70]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[306]}), .b4_nUAi({
        b4_nUAi[212], b4_nUAi[211], b4_nUAi[210]}), .b6_2ZTGIf({
        \b6_2ZTGIf[70] }));
    b8_1LbcQDr1_x_366_0 b8_1LbcgKGR (.mdiclink_reg({mdiclink_reg[10]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[366]}), .b4_nUAi({
        b4_nUAi[32], b4_nUAi[31], b4_nUAi[30]}), .b6_2ZTGIf({
        \b6_2ZTGIf[10] }));
    b8_1LbcQDr1_x_204_0 b9_1LbcgKGJd (.mdiclink_reg({mdiclink_reg[172]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[204]}), .b4_nUAi({
        b4_nUAi[517], b4_nUAi[516]}), .N_27(N_27_61), .N_25(N_25_61));
    b8_1LbcQDr1_x_325_0 b8_1LbcgKIS (.mdiclink_reg({mdiclink_reg[51]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[325]}), .b4_nUAi({
        b4_nUAi[155], b4_nUAi[154], b4_nUAi[153]}), .b6_2ZTGIf({
        \b6_2ZTGIf[51] }));
    b16_CRGcTCua_eH4_2j7_x_0 b6_2ZGFQ9 (.b11_uUT0JC4gFrY({
        b11_uUT0JC4gFrY[1]}), .b4_nUAi_0(b4_nUAi[17]), .b4_nUAi_30(
        b4_nUAi[47]), .b4_nUAi_27(b4_nUAi[44]), .b4_nUAi_24(
        b4_nUAi[41]), .b4_nUAi_21(b4_nUAi[38]), .b4_nUAi_18(
        b4_nUAi[35]), .b4_nUAi_48(b4_nUAi[65]), .b4_nUAi_78(
        b4_nUAi[95]), .b4_nUAi_75(b4_nUAi[92]), .b4_nUAi_72(
        b4_nUAi[89]), .b4_nUAi_69(b4_nUAi[86]), .b4_nUAi_66(
        b4_nUAi[83]), .b4_nUAi_96(b4_nUAi[113]), .b4_nUAi_126(
        b4_nUAi[143]), .b4_nUAi_123(b4_nUAi[140]), .b4_nUAi_120(
        b4_nUAi[137]), .b4_nUAi_117(b4_nUAi[134]), .b4_nUAi_114(
        b4_nUAi[131]), .b4_nUAi_144(b4_nUAi[161]), .b4_nUAi_174(
        b4_nUAi[191]), .b4_nUAi_171(b4_nUAi[188]), .b4_nUAi_168(
        b4_nUAi[185]), .b4_nUAi_165(b4_nUAi[182]), .b4_nUAi_162(
        b4_nUAi[179]), .b4_nUAi_192(b4_nUAi[209]), .b4_nUAi_222(
        b4_nUAi[239]), .b4_nUAi_219(b4_nUAi[236]), .b4_nUAi_216(
        b4_nUAi[233]), .b4_nUAi_213(b4_nUAi[230]), .b4_nUAi_210(
        b4_nUAi[227]), .b4_nUAi_240(b4_nUAi[257]), .b4_nUAi_270(
        b4_nUAi[287]), .b4_nUAi_267(b4_nUAi[284]), .b4_nUAi_264(
        b4_nUAi[281]), .b4_nUAi_261(b4_nUAi[278]), .b4_nUAi_258(
        b4_nUAi[275]), .b4_nUAi_288(b4_nUAi[305]), .b4_nUAi_318(
        b4_nUAi[335]), .b4_nUAi_315(b4_nUAi[332]), .b4_nUAi_312(
        b4_nUAi[329]), .b4_nUAi_309(b4_nUAi[326]), .b4_nUAi_306(
        b4_nUAi[323]), .b4_nUAi_336(b4_nUAi[353]), .b4_nUAi_366(
        b4_nUAi[383]), .b4_nUAi_363(b4_nUAi[380]), .b4_nUAi_360(
        b4_nUAi[377]), .b4_nUAi_357(b4_nUAi[374]), .b4_nUAi_354(
        b4_nUAi[371]), .b4_nUAi_384(b4_nUAi[401]), .b4_nUAi_414(
        b4_nUAi[431]), .b4_nUAi_411(b4_nUAi[428]), .b4_nUAi_408(
        b4_nUAi[425]), .b4_nUAi_405(b4_nUAi[422]), .b4_nUAi_402(
        b4_nUAi[419]), .b4_nUAi_432(b4_nUAi[449]), .b4_nUAi_462(
        b4_nUAi[479]), .b4_nUAi_459(b4_nUAi[476]), .b4_nUAi_456(
        b4_nUAi[473]), .b4_nUAi_453(b4_nUAi[470]), .b4_nUAi_450(
        b4_nUAi[467]), .b4_nUAi_480(b4_nUAi[497]), .b4_nUAi_510(
        b4_nUAi[527]), .b4_nUAi_507(b4_nUAi[524]), .b4_nUAi_504(
        b4_nUAi[521]), .b4_nUAi_501(b4_nUAi[518]), .b4_nUAi_498(
        b4_nUAi[515]), .b4_nUAi_528(b4_nUAi[545]), .b4_nUAi_558(
        b4_nUAi[575]), .b4_nUAi_555(b4_nUAi[572]), .b4_nUAi_552(
        b4_nUAi[569]), .b4_nUAi_549(b4_nUAi[566]), .b4_nUAi_546(
        b4_nUAi[563]), .b4_nUAi_576(b4_nUAi[593]), .b4_nUAi_606(
        b4_nUAi[623]), .b4_nUAi_603(b4_nUAi[620]), .b4_nUAi_600(
        b4_nUAi[617]), .b4_nUAi_597(b4_nUAi[614]), .b4_nUAi_594(
        b4_nUAi[611]), .b4_nUAi_624(b4_nUAi[641]), .b4_nUAi_654(
        b4_nUAi[671]), .b4_nUAi_651(b4_nUAi[668]), .b4_nUAi_648(
        b4_nUAi[665]), .b4_nUAi_645(b4_nUAi[662]), .b4_nUAi_642(
        b4_nUAi[659]), .b4_nUAi_672(b4_nUAi[689]), .b4_nUAi_702(
        b4_nUAi[719]), .b4_nUAi_699(b4_nUAi[716]), .b4_nUAi_696(
        b4_nUAi[713]), .b4_nUAi_693(b4_nUAi[710]), .b4_nUAi_690(
        b4_nUAi[707]), .b4_nUAi_720(b4_nUAi[737]), .b4_nUAi_750(
        b4_nUAi[767]), .b4_nUAi_747(b4_nUAi[764]), .b4_nUAi_744(
        b4_nUAi[761]), .b4_nUAi_741(b4_nUAi[758]), .b4_nUAi_738(
        b4_nUAi[755]), .b4_nUAi_768(b4_nUAi[785]), .b4_nUAi_798(
        b4_nUAi[815]), .b4_nUAi_795(b4_nUAi[812]), .b4_nUAi_792(
        b4_nUAi[809]), .b4_nUAi_789(b4_nUAi[806]), .b4_nUAi_786(
        b4_nUAi[803]), .b4_nUAi_816(b4_nUAi[833]), .b4_nUAi_846(
        b4_nUAi[863]), .b4_nUAi_843(b4_nUAi[860]), .b4_nUAi_840(
        b4_nUAi[857]), .b4_nUAi_837(b4_nUAi[854]), .b4_nUAi_834(
        b4_nUAi[851]), .b4_nUAi_864(b4_nUAi[881]), .b4_nUAi_894(
        b4_nUAi[911]), .b4_nUAi_891(b4_nUAi[908]), .b4_nUAi_888(
        b4_nUAi[905]), .b4_nUAi_885(b4_nUAi[902]), .b4_nUAi_882(
        b4_nUAi[899]), .b4_nUAi_912(b4_nUAi[929]), .b4_nUAi_942(
        b4_nUAi[959]), .b4_nUAi_939(b4_nUAi[956]), .b4_nUAi_936(
        b4_nUAi[953]), .b4_nUAi_933(b4_nUAi[950]), .b4_nUAi_930(
        b4_nUAi[947]), .b4_nUAi_960(b4_nUAi[977]), .b4_nUAi_990(
        b4_nUAi[1007]), .b4_nUAi_987(b4_nUAi[1004]), .b4_nUAi_984(
        b4_nUAi[1001]), .b4_nUAi_981(b4_nUAi[998]), .b4_nUAi_978(
        b4_nUAi[995]), .b4_nUAi_1008(b4_nUAi[1025]), .b4_nUAi_1038(
        b4_nUAi[1055]), .b4_nUAi_1035(b4_nUAi[1052]), .b4_nUAi_1032(
        b4_nUAi[1049]), .b4_nUAi_1029(b4_nUAi[1046]), .b4_nUAi_1026(
        b4_nUAi[1043]), .b4_nUAi_1056(b4_nUAi[1073]), .b4_nUAi_1086(
        b4_nUAi[1103]), .b4_nUAi_1083(b4_nUAi[1100]), .b4_nUAi_1080(
        b4_nUAi[1097]), .b4_nUAi_1077(b4_nUAi[1094]), .b4_nUAi_1074(
        b4_nUAi[1091]), .b4_nUAi_1107(b4_nUAi[1124]), .b4_nUAi_1101(
        b4_nUAi[1118]), .b4_nUAi_1095(b4_nUAi[1112]), .b4_nUAi_1089(
        b4_nUAi[1106]), .b6_2ZTGIf_6(\b6_2ZTGIf[6] ), .b6_2ZTGIf_4(
        \b6_2ZTGIf[4] ), .b6_2ZTGIf_3(\b6_2ZTGIf[3] ), .b6_2ZTGIf_2(
        \b6_2ZTGIf[2] ), .b6_2ZTGIf_1(\b6_2ZTGIf[1] ), .b6_2ZTGIf_0(
        \b6_2ZTGIf[0] ), .b6_2ZTGIf_10(\b6_2ZTGIf[10] ), .b6_2ZTGIf_9(
        \b6_2ZTGIf[9] ), .b6_2ZTGIf_8(\b6_2ZTGIf[8] ), .b6_2ZTGIf_7(
        \b6_2ZTGIf[7] ), .b6_2ZTGIf_22(\b6_2ZTGIf[22] ), .b6_2ZTGIf_20(
        \b6_2ZTGIf[20] ), .b6_2ZTGIf_19(\b6_2ZTGIf[19] ), 
        .b6_2ZTGIf_18(\b6_2ZTGIf[18] ), .b6_2ZTGIf_17(\b6_2ZTGIf[17] ), 
        .b6_2ZTGIf_16(\b6_2ZTGIf[16] ), .b6_2ZTGIf_26(\b6_2ZTGIf[26] ), 
        .b6_2ZTGIf_25(\b6_2ZTGIf[25] ), .b6_2ZTGIf_24(\b6_2ZTGIf[24] ), 
        .b6_2ZTGIf_23(\b6_2ZTGIf[23] ), .b6_2ZTGIf_38(\b6_2ZTGIf[38] ), 
        .b6_2ZTGIf_36(\b6_2ZTGIf[36] ), .b6_2ZTGIf_35(\b6_2ZTGIf[35] ), 
        .b6_2ZTGIf_34(\b6_2ZTGIf[34] ), .b6_2ZTGIf_33(\b6_2ZTGIf[33] ), 
        .b6_2ZTGIf_32(\b6_2ZTGIf[32] ), .b6_2ZTGIf_42(\b6_2ZTGIf[42] ), 
        .b6_2ZTGIf_41(\b6_2ZTGIf[41] ), .b6_2ZTGIf_40(\b6_2ZTGIf[40] ), 
        .b6_2ZTGIf_39(\b6_2ZTGIf[39] ), .b6_2ZTGIf_54(\b6_2ZTGIf[54] ), 
        .b6_2ZTGIf_52(\b6_2ZTGIf[52] ), .b6_2ZTGIf_51(\b6_2ZTGIf[51] ), 
        .b6_2ZTGIf_50(\b6_2ZTGIf[50] ), .b6_2ZTGIf_49(\b6_2ZTGIf[49] ), 
        .b6_2ZTGIf_48(\b6_2ZTGIf[48] ), .b6_2ZTGIf_58(\b6_2ZTGIf[58] ), 
        .b6_2ZTGIf_57(\b6_2ZTGIf[57] ), .b6_2ZTGIf_56(\b6_2ZTGIf[56] ), 
        .b6_2ZTGIf_55(\b6_2ZTGIf[55] ), .b6_2ZTGIf_70(\b6_2ZTGIf[70] ), 
        .b6_2ZTGIf_68(\b6_2ZTGIf[68] ), .b6_2ZTGIf_67(\b6_2ZTGIf[67] ), 
        .b6_2ZTGIf_66(\b6_2ZTGIf[66] ), .b6_2ZTGIf_65(\b6_2ZTGIf[65] ), 
        .b6_2ZTGIf_64(\b6_2ZTGIf[64] ), .b6_2ZTGIf_74(\b6_2ZTGIf[74] ), 
        .b6_2ZTGIf_73(\b6_2ZTGIf[73] ), .b6_2ZTGIf_72(\b6_2ZTGIf[72] ), 
        .b6_2ZTGIf_71(\b6_2ZTGIf[71] ), .b6_2ZTGIf_86(\b6_2ZTGIf[86] ), 
        .b6_2ZTGIf_84(\b6_2ZTGIf[84] ), .b6_2ZTGIf_83(\b6_2ZTGIf[83] ), 
        .b6_2ZTGIf_82(\b6_2ZTGIf[82] ), .b6_2ZTGIf_81(\b6_2ZTGIf[81] ), 
        .b6_2ZTGIf_80(\b6_2ZTGIf[80] ), .b6_2ZTGIf_90(\b6_2ZTGIf[90] ), 
        .b6_2ZTGIf_89(\b6_2ZTGIf[89] ), .b6_2ZTGIf_88(\b6_2ZTGIf[88] ), 
        .b6_2ZTGIf_87(\b6_2ZTGIf[87] ), .b6_2ZTGIf_102(
        \b6_2ZTGIf[102] ), .b6_2ZTGIf_100(\b6_2ZTGIf[100] ), 
        .b6_2ZTGIf_99(\b6_2ZTGIf[99] ), .b6_2ZTGIf_98(\b6_2ZTGIf[98] ), 
        .b6_2ZTGIf_97(\b6_2ZTGIf[97] ), .b6_2ZTGIf_96(\b6_2ZTGIf[96] ), 
        .b6_2ZTGIf_106(\b6_2ZTGIf[106] ), .b6_2ZTGIf_105(
        \b6_2ZTGIf[105] ), .b6_2ZTGIf_104(\b6_2ZTGIf[104] ), 
        .b6_2ZTGIf_103(\b6_2ZTGIf[103] ), .b6_2ZTGIf_118(
        \b6_2ZTGIf[118] ), .b6_2ZTGIf_116(\b6_2ZTGIf[116] ), 
        .b6_2ZTGIf_115(\b6_2ZTGIf[115] ), .b6_2ZTGIf_114(
        \b6_2ZTGIf[114] ), .b6_2ZTGIf_113(\b6_2ZTGIf[113] ), 
        .b6_2ZTGIf_112(\b6_2ZTGIf[112] ), .b6_2ZTGIf_122(
        \b6_2ZTGIf[122] ), .b6_2ZTGIf_121(\b6_2ZTGIf[121] ), 
        .b6_2ZTGIf_120(\b6_2ZTGIf[120] ), .b6_2ZTGIf_119(
        \b6_2ZTGIf[119] ), .b6_2ZTGIf_134(\b6_2ZTGIf[134] ), 
        .b6_2ZTGIf_132(\b6_2ZTGIf[132] ), .b6_2ZTGIf_131(
        \b6_2ZTGIf[131] ), .b6_2ZTGIf_130(\b6_2ZTGIf[130] ), 
        .b6_2ZTGIf_129(\b6_2ZTGIf[129] ), .b6_2ZTGIf_128(
        \b6_2ZTGIf[128] ), .b6_2ZTGIf_138(\b6_2ZTGIf[138] ), 
        .b6_2ZTGIf_137(\b6_2ZTGIf[137] ), .b6_2ZTGIf_136(
        \b6_2ZTGIf[136] ), .b6_2ZTGIf_135(\b6_2ZTGIf[135] ), 
        .b6_2ZTGIf_150(\b6_2ZTGIf[150] ), .b6_2ZTGIf_148(
        \b6_2ZTGIf[148] ), .b6_2ZTGIf_147(\b6_2ZTGIf[147] ), 
        .b6_2ZTGIf_146(\b6_2ZTGIf[146] ), .b6_2ZTGIf_145(
        \b6_2ZTGIf[145] ), .b6_2ZTGIf_144(\b6_2ZTGIf[144] ), 
        .b6_2ZTGIf_154(\b6_2ZTGIf[154] ), .b6_2ZTGIf_153(
        \b6_2ZTGIf[153] ), .b6_2ZTGIf_152(\b6_2ZTGIf[152] ), 
        .b6_2ZTGIf_151(\b6_2ZTGIf[151] ), .b6_2ZTGIf_166(
        \b6_2ZTGIf[166] ), .b6_2ZTGIf_164(\b6_2ZTGIf[164] ), 
        .b6_2ZTGIf_163(\b6_2ZTGIf[163] ), .b6_2ZTGIf_162(
        \b6_2ZTGIf[162] ), .b6_2ZTGIf_161(\b6_2ZTGIf[161] ), 
        .b6_2ZTGIf_160(\b6_2ZTGIf[160] ), .b6_2ZTGIf_170(
        \b6_2ZTGIf[170] ), .b6_2ZTGIf_169(\b6_2ZTGIf[169] ), 
        .b6_2ZTGIf_168(\b6_2ZTGIf[168] ), .b6_2ZTGIf_167(
        \b6_2ZTGIf[167] ), .b6_2ZTGIf_182(\b6_2ZTGIf[182] ), 
        .b6_2ZTGIf_180(\b6_2ZTGIf[180] ), .b6_2ZTGIf_179(
        \b6_2ZTGIf[179] ), .b6_2ZTGIf_178(\b6_2ZTGIf[178] ), 
        .b6_2ZTGIf_177(\b6_2ZTGIf[177] ), .b6_2ZTGIf_176(
        \b6_2ZTGIf[176] ), .b6_2ZTGIf_186(\b6_2ZTGIf[186] ), 
        .b6_2ZTGIf_185(\b6_2ZTGIf[185] ), .b6_2ZTGIf_184(
        \b6_2ZTGIf[184] ), .b6_2ZTGIf_183(\b6_2ZTGIf[183] ), 
        .b6_2ZTGIf_198(\b6_2ZTGIf[198] ), .b6_2ZTGIf_196(
        \b6_2ZTGIf[196] ), .b6_2ZTGIf_195(\b6_2ZTGIf[195] ), 
        .b6_2ZTGIf_194(\b6_2ZTGIf[194] ), .b6_2ZTGIf_193(
        \b6_2ZTGIf[193] ), .b6_2ZTGIf_192(\b6_2ZTGIf[192] ), 
        .b6_2ZTGIf_202(\b6_2ZTGIf[202] ), .b6_2ZTGIf_201(
        \b6_2ZTGIf[201] ), .b6_2ZTGIf_200(\b6_2ZTGIf[200] ), 
        .b6_2ZTGIf_199(\b6_2ZTGIf[199] ), .b6_2ZTGIf_214(
        \b6_2ZTGIf[214] ), .b6_2ZTGIf_212(\b6_2ZTGIf[212] ), 
        .b6_2ZTGIf_211(\b6_2ZTGIf[211] ), .b6_2ZTGIf_210(
        \b6_2ZTGIf[210] ), .b6_2ZTGIf_209(\b6_2ZTGIf[209] ), 
        .b6_2ZTGIf_208(\b6_2ZTGIf[208] ), .b6_2ZTGIf_218(
        \b6_2ZTGIf[218] ), .b6_2ZTGIf_217(\b6_2ZTGIf[217] ), 
        .b6_2ZTGIf_216(\b6_2ZTGIf[216] ), .b6_2ZTGIf_215(
        \b6_2ZTGIf[215] ), .b6_2ZTGIf_230(\b6_2ZTGIf[230] ), 
        .b6_2ZTGIf_228(\b6_2ZTGIf[228] ), .b6_2ZTGIf_227(
        \b6_2ZTGIf[227] ), .b6_2ZTGIf_226(\b6_2ZTGIf[226] ), 
        .b6_2ZTGIf_225(\b6_2ZTGIf[225] ), .b6_2ZTGIf_224(
        \b6_2ZTGIf[224] ), .b6_2ZTGIf_234(\b6_2ZTGIf[234] ), 
        .b6_2ZTGIf_233(\b6_2ZTGIf[233] ), .b6_2ZTGIf_232(
        \b6_2ZTGIf[232] ), .b6_2ZTGIf_231(\b6_2ZTGIf[231] ), 
        .b6_2ZTGIf_246(\b6_2ZTGIf[246] ), .b6_2ZTGIf_244(
        \b6_2ZTGIf[244] ), .b6_2ZTGIf_243(\b6_2ZTGIf[243] ), 
        .b6_2ZTGIf_242(\b6_2ZTGIf[242] ), .b6_2ZTGIf_241(
        \b6_2ZTGIf[241] ), .b6_2ZTGIf_240(\b6_2ZTGIf[240] ), 
        .b6_2ZTGIf_250(\b6_2ZTGIf[250] ), .b6_2ZTGIf_249(
        \b6_2ZTGIf[249] ), .b6_2ZTGIf_248(\b6_2ZTGIf[248] ), 
        .b6_2ZTGIf_247(\b6_2ZTGIf[247] ), .b6_2ZTGIf_262(
        \b6_2ZTGIf[262] ), .b6_2ZTGIf_260(\b6_2ZTGIf[260] ), 
        .b6_2ZTGIf_259(\b6_2ZTGIf[259] ), .b6_2ZTGIf_258(
        \b6_2ZTGIf[258] ), .b6_2ZTGIf_257(\b6_2ZTGIf[257] ), 
        .b6_2ZTGIf_256(\b6_2ZTGIf[256] ), .b6_2ZTGIf_266(
        \b6_2ZTGIf[266] ), .b6_2ZTGIf_265(\b6_2ZTGIf[265] ), 
        .b6_2ZTGIf_264(\b6_2ZTGIf[264] ), .b6_2ZTGIf_263(
        \b6_2ZTGIf[263] ), .b6_2ZTGIf_278(\b6_2ZTGIf[278] ), 
        .b6_2ZTGIf_276(\b6_2ZTGIf[276] ), .b6_2ZTGIf_275(
        \b6_2ZTGIf[275] ), .b6_2ZTGIf_274(\b6_2ZTGIf[274] ), 
        .b6_2ZTGIf_273(\b6_2ZTGIf[273] ), .b6_2ZTGIf_272(
        \b6_2ZTGIf[272] ), .b6_2ZTGIf_282(\b6_2ZTGIf[282] ), 
        .b6_2ZTGIf_281(\b6_2ZTGIf[281] ), .b6_2ZTGIf_280(
        \b6_2ZTGIf[280] ), .b6_2ZTGIf_279(\b6_2ZTGIf[279] ), 
        .b6_2ZTGIf_294(\b6_2ZTGIf[294] ), .b6_2ZTGIf_292(
        \b6_2ZTGIf[292] ), .b6_2ZTGIf_291(\b6_2ZTGIf[291] ), 
        .b6_2ZTGIf_290(\b6_2ZTGIf[290] ), .b6_2ZTGIf_289(
        \b6_2ZTGIf[289] ), .b6_2ZTGIf_288(\b6_2ZTGIf[288] ), 
        .b6_2ZTGIf_298(\b6_2ZTGIf[298] ), .b6_2ZTGIf_297(
        \b6_2ZTGIf[297] ), .b6_2ZTGIf_296(\b6_2ZTGIf[296] ), 
        .b6_2ZTGIf_295(\b6_2ZTGIf[295] ), .b6_2ZTGIf_310(
        \b6_2ZTGIf[310] ), .b6_2ZTGIf_308(\b6_2ZTGIf[308] ), 
        .b6_2ZTGIf_307(\b6_2ZTGIf[307] ), .b6_2ZTGIf_306(
        \b6_2ZTGIf[306] ), .b6_2ZTGIf_305(\b6_2ZTGIf[305] ), 
        .b6_2ZTGIf_304(\b6_2ZTGIf[304] ), .b6_2ZTGIf_314(
        \b6_2ZTGIf[314] ), .b6_2ZTGIf_313(\b6_2ZTGIf[313] ), 
        .b6_2ZTGIf_312(\b6_2ZTGIf[312] ), .b6_2ZTGIf_311(
        \b6_2ZTGIf[311] ), .b6_2ZTGIf_326(\b6_2ZTGIf[326] ), 
        .b6_2ZTGIf_324(\b6_2ZTGIf[324] ), .b6_2ZTGIf_323(
        \b6_2ZTGIf[323] ), .b6_2ZTGIf_322(\b6_2ZTGIf[322] ), 
        .b6_2ZTGIf_321(\b6_2ZTGIf[321] ), .b6_2ZTGIf_320(
        \b6_2ZTGIf[320] ), .b6_2ZTGIf_330(\b6_2ZTGIf[330] ), 
        .b6_2ZTGIf_329(\b6_2ZTGIf[329] ), .b6_2ZTGIf_328(
        \b6_2ZTGIf[328] ), .b6_2ZTGIf_327(\b6_2ZTGIf[327] ), 
        .b6_2ZTGIf_342(\b6_2ZTGIf[342] ), .b6_2ZTGIf_340(
        \b6_2ZTGIf[340] ), .b6_2ZTGIf_339(\b6_2ZTGIf[339] ), 
        .b6_2ZTGIf_338(\b6_2ZTGIf[338] ), .b6_2ZTGIf_337(
        \b6_2ZTGIf[337] ), .b6_2ZTGIf_336(\b6_2ZTGIf[336] ), 
        .b6_2ZTGIf_346(\b6_2ZTGIf[346] ), .b6_2ZTGIf_345(
        \b6_2ZTGIf[345] ), .b6_2ZTGIf_344(\b6_2ZTGIf[344] ), 
        .b6_2ZTGIf_343(\b6_2ZTGIf[343] ), .b6_2ZTGIf_358(
        \b6_2ZTGIf[358] ), .b6_2ZTGIf_356(\b6_2ZTGIf[356] ), 
        .b6_2ZTGIf_355(\b6_2ZTGIf[355] ), .b6_2ZTGIf_354(
        \b6_2ZTGIf[354] ), .b6_2ZTGIf_353(\b6_2ZTGIf[353] ), 
        .b6_2ZTGIf_352(\b6_2ZTGIf[352] ), .b6_2ZTGIf_362(
        \b6_2ZTGIf[362] ), .b6_2ZTGIf_361(\b6_2ZTGIf[361] ), 
        .b6_2ZTGIf_360(\b6_2ZTGIf[360] ), .b6_2ZTGIf_359(
        \b6_2ZTGIf[359] ), .b6_2ZTGIf_375(\b6_2ZTGIf[375] ), 
        .b6_2ZTGIf_373(\b6_2ZTGIf[373] ), .b6_2ZTGIf_371(
        \b6_2ZTGIf[371] ), .b6_2ZTGIf_369(\b6_2ZTGIf[369] ), .BW_clk_c(
        BW_clk_c), .N_25(N_25), .N_27(N_27), .N_25_0(N_25_4), .N_27_0(
        N_27_4), .N_25_1(N_25_3), .N_27_1(N_27_3), .N_25_2(N_25_2), 
        .N_27_2(N_27_2), .N_25_3(N_25_1), .N_27_3(N_27_1), .N_25_4(
        N_25_0), .N_27_4(N_27_0), .N_25_5(N_25_5), .N_27_5(N_27_5), 
        .N_25_6(N_25_10), .N_27_6(N_27_10), .N_25_7(N_25_9), .N_27_7(
        N_27_9), .N_25_8(N_25_8), .N_27_8(N_27_8), .N_25_9(N_25_7), 
        .N_27_9(N_27_7), .N_25_10(N_25_6), .N_27_10(N_27_6), .N_25_11(
        N_25_11), .N_27_11(N_27_11), .N_25_12(N_25_16), .N_27_12(
        N_27_16), .N_25_13(N_25_15), .N_27_13(N_27_15), .N_25_14(
        N_25_14), .N_27_14(N_27_14), .N_25_15(N_25_13), .N_27_15(
        N_27_13), .N_25_16(N_25_12), .N_27_16(N_27_12), .N_25_17(
        N_25_17), .N_27_17(N_27_17), .N_25_18(N_25_22), .N_27_18(
        N_27_22), .N_25_19(N_25_21), .N_27_19(N_27_21), .N_25_20(
        N_25_20), .N_27_20(N_27_20), .N_25_21(N_25_19), .N_27_21(
        N_27_19), .N_25_22(N_25_18), .N_27_22(N_27_18), .N_25_23(
        N_25_23), .N_27_23(N_27_23), .N_25_24(N_25_28), .N_27_24(
        N_27_28), .N_25_25(N_25_27), .N_27_25(N_27_27), .N_25_26(
        N_25_26), .N_27_26(N_27_26), .N_25_27(N_25_25), .N_27_27(
        N_27_25), .N_25_28(N_25_24), .N_27_28(N_27_24), .N_25_29(
        N_25_29), .N_27_29(N_27_29), .N_25_30(N_25_34), .N_27_30(
        N_27_34), .N_25_31(N_25_33), .N_27_31(N_27_33), .N_25_32(
        N_25_32), .N_27_32(N_27_32), .N_25_33(N_25_31), .N_27_33(
        N_27_31), .N_25_34(N_25_30), .N_27_34(N_27_30), .N_25_35(
        N_25_35), .N_27_35(N_27_35), .N_25_36(N_25_40), .N_27_36(
        N_27_40), .N_25_37(N_25_39), .N_27_37(N_27_39), .N_25_38(
        N_25_38), .N_27_38(N_27_38), .N_25_39(N_25_37), .N_27_39(
        N_27_37), .N_25_40(N_25_36), .N_27_40(N_27_36), .N_25_41(
        N_25_41), .N_27_41(N_27_41), .N_25_42(N_25_46), .N_27_42(
        N_27_46), .N_25_43(N_25_45), .N_27_43(N_27_45), .N_25_44(
        N_25_44), .N_27_44(N_27_44), .N_25_45(N_25_43), .N_27_45(
        N_27_43), .N_25_46(N_25_42), .N_27_46(N_27_42), .N_25_47(
        N_25_47), .N_27_47(N_27_47), .N_25_48(N_25_52), .N_27_48(
        N_27_52), .N_25_49(N_25_51), .N_27_49(N_27_51), .N_25_50(
        N_25_50), .N_27_50(N_27_50), .N_25_51(N_25_49), .N_27_51(
        N_27_49), .N_25_52(N_25_48), .N_27_52(N_27_48), .N_25_53(
        N_25_53), .N_27_53(N_27_53), .N_25_54(N_25_58), .N_27_54(
        N_27_58), .N_25_55(N_25_57), .N_27_55(N_27_57), .N_25_56(
        N_25_56), .N_27_56(N_27_56), .N_25_57(N_25_55), .N_27_57(
        N_27_55), .N_25_58(N_25_54), .N_27_58(N_27_54), .N_25_59(
        N_25_59), .N_27_59(N_27_59), .N_25_60(N_25_64), .N_27_60(
        N_27_64), .N_25_61(N_25_63), .N_27_61(N_27_63), .N_25_62(
        N_25_62), .N_27_62(N_27_62), .N_25_63(N_25_61), .N_27_63(
        N_27_61), .N_25_64(N_25_60), .N_27_64(N_27_60), .N_25_65(
        N_25_65), .N_27_65(N_27_65), .N_25_66(N_25_70), .N_27_66(
        N_27_70), .N_25_67(N_25_69), .N_27_67(N_27_69), .N_25_68(
        N_25_68), .N_27_68(N_27_68), .N_25_69(N_25_67), .N_27_69(
        N_27_67), .N_25_70(N_25_66), .N_27_70(N_27_66), .N_25_71(
        N_25_71), .N_27_71(N_27_71), .N_25_72(N_25_76), .N_27_72(
        N_27_76), .N_25_73(N_25_75), .N_27_73(N_27_75), .N_25_74(
        N_25_74), .N_27_74(N_27_74), .N_25_75(N_25_73), .N_27_75(
        N_27_73), .N_25_76(N_25_72), .N_27_76(N_27_72), .N_25_77(
        N_25_77), .N_27_77(N_27_77), .N_25_78(N_25_82), .N_27_78(
        N_27_82), .N_25_79(N_25_81), .N_27_79(N_27_81), .N_25_80(
        N_25_80), .N_27_80(N_27_80), .N_25_81(N_25_79), .N_27_81(
        N_27_79), .N_25_82(N_25_78), .N_27_82(N_27_78), .N_25_83(
        N_25_83), .N_27_83(N_27_83), .N_25_84(N_25_88), .N_27_84(
        N_27_88), .N_25_85(N_25_87), .N_27_85(N_27_87), .N_25_86(
        N_25_86), .N_27_86(N_27_86), .N_25_87(N_25_85), .N_27_87(
        N_27_85), .N_25_88(N_25_84), .N_27_88(N_27_84), .N_25_89(
        N_25_89), .N_27_89(N_27_89), .N_25_90(N_25_94), .N_27_90(
        N_27_94), .N_25_91(N_25_93), .N_27_91(N_27_93), .N_25_92(
        N_25_92), .N_27_92(N_27_92), .N_25_93(N_25_91), .N_27_93(
        N_27_91), .N_25_94(N_25_90), .N_27_94(N_27_90), .N_25_95(
        N_25_95), .N_27_95(N_27_95), .N_25_96(N_25_100), .N_27_96(
        N_27_100), .N_25_97(N_25_99), .N_27_97(N_27_99), .N_25_98(
        N_25_98), .N_27_98(N_27_98), .N_25_99(N_25_97), .N_27_99(
        N_27_97), .N_25_100(N_25_96), .N_27_100(N_27_96), .N_25_101(
        N_25_101), .N_27_101(N_27_101), .N_25_102(N_25_106), .N_27_102(
        N_27_106), .N_25_103(N_25_105), .N_27_103(N_27_105), .N_25_104(
        N_25_104), .N_27_104(N_27_104), .N_25_105(N_25_103), .N_27_105(
        N_27_103), .N_25_106(N_25_102), .N_27_106(N_27_102), .N_25_107(
        N_25_107), .N_27_107(N_27_107), .N_25_108(N_25_112), .N_27_108(
        N_27_112), .N_25_109(N_25_111), .N_27_109(N_27_111), .N_25_110(
        N_25_110), .N_27_110(N_27_110), .N_25_111(N_25_109), .N_27_111(
        N_27_109), .N_25_112(N_25_108), .N_27_112(N_27_108), .N_25_113(
        N_25_113), .N_27_113(N_27_113), .N_25_114(N_25_118), .N_27_114(
        N_27_118), .N_25_115(N_25_117), .N_27_115(N_27_117), .N_25_116(
        N_25_116), .N_27_116(N_27_116), .N_25_117(N_25_115), .N_27_117(
        N_27_115), .N_25_118(N_25_114), .N_27_118(N_27_114), .N_25_119(
        N_25_119), .N_27_119(N_27_119), .N_25_120(N_25_124), .N_27_120(
        N_27_124), .N_25_121(N_25_123), .N_27_121(N_27_123), .N_25_122(
        N_25_122), .N_27_122(N_27_122), .N_25_123(N_25_121), .N_27_123(
        N_27_121), .N_25_124(N_25_120), .N_27_124(N_27_120), .N_25_125(
        N_25_125), .N_27_125(N_27_125), .N_25_126(N_25_130), .N_27_126(
        N_27_130), .N_25_127(N_25_129), .N_27_127(N_27_129), .N_25_128(
        N_25_128), .N_27_128(N_27_128), .N_25_129(N_25_127), .N_27_129(
        N_27_127), .N_25_130(N_25_126), .N_27_130(N_27_126), .N_25_131(
        N_25_131), .N_27_131(N_27_131), .N_25_132(N_25_136), .N_27_132(
        N_27_136), .N_25_133(N_25_135), .N_27_133(N_27_135), .N_25_134(
        N_25_134), .N_27_134(N_27_134), .N_25_135(N_25_133), .N_27_135(
        N_27_133), .N_25_136(N_25_132), .N_27_136(N_27_132), .N_25_137(
        N_25_140), .N_27_137(N_27_140), .N_25_138(N_25_139), .N_27_138(
        N_27_139), .N_25_139(N_25_138), .N_27_139(N_27_138), .N_25_140(
        N_25_137), .N_27_140(N_27_137), .N_25_141(N_25_141), 
        .b7_PSyi3wy(b7_PSyi3wy), .N_27_141(N_27_141));
    b8_1LbcQDr1_x_51_0 b9_1LbcgKeIp (.mdiclink_reg({mdiclink_reg[325]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[51]}), .b4_nUAi({
        b4_nUAi[976], b4_nUAi[975]}), .N_27(N_27_119), .N_25(N_25_119));
    b8_1LbcQDr1_x_326_0 b8_1LbcgKIR (.mdiclink_reg({mdiclink_reg[50]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[326]}), .b4_nUAi({
        b4_nUAi[152], b4_nUAi[151], b4_nUAi[150]}), .b6_2ZTGIf({
        \b6_2ZTGIf[50] }));
    b8_1LbcQDr1_x_294_0 b8_1LbcgKbI (.mdiclink_reg({mdiclink_reg[82]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[294]}), .b4_nUAi({
        b4_nUAi[248], b4_nUAi[247], b4_nUAi[246]}), .b6_2ZTGIf({
        \b6_2ZTGIf[82] }));
    b8_1LbcQDr1_x_8_0 b9_1LbcgKeAS (.mdiclink_reg({mdiclink_reg[368]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[8]}), .b4_nUAi({
        b4_nUAi[1105], b4_nUAi[1104]}), .N_27(N_27_137), .N_25(
        N_25_137));
    b8_1LbcQDr1_x_65_0 b9_1LbcgKeSn (.mdiclink_reg({mdiclink_reg[311]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[65]}), .b4_nUAi({
        b4_nUAi[935], b4_nUAi[934], b4_nUAi[933]}), .b6_2ZTGIf({
        \b6_2ZTGIf[311] }));
    b8_1LbcQDr1_x_75_0 b9_1LbcgKeRn (.mdiclink_reg({mdiclink_reg[301]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[75]}), .b4_nUAi({
        b4_nUAi[904], b4_nUAi[903]}), .N_27(N_27_110), .N_25(N_25_110));
    b8_1LbcQDr1_x_138_0 b9_1LbcgKwqS (.mdiclink_reg({mdiclink_reg[238]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[138]}), .b4_nUAi({
        b4_nUAi[715], b4_nUAi[714]}), .N_27(N_27_87), .N_25(N_25_87));
    b8_1LbcQDr1_x_255_0 b9_1LbcgKGIn (.mdiclink_reg({mdiclink_reg[121]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[255]}), .b4_nUAi({
        b4_nUAi[365], b4_nUAi[364], b4_nUAi[363]}), .b6_2ZTGIf({
        \b6_2ZTGIf[121] }));
    b8_1LbcQDr1_x_92_0 b9_1LbcgKwnl (.mdiclink_reg({mdiclink_reg[284]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[92]}), .b4_nUAi({
        b4_nUAi[853], b4_nUAi[852]}), .N_27(N_27_103), .N_25(N_25_103));
    b8_1LbcQDr1_x_28_0 b9_1LbcgKeQS0 (.mdiclink_reg({mdiclink_reg[348]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[28]}), .b4_nUAi({
        b4_nUAi[1045], b4_nUAi[1044]}), .N_27(N_27_127), .N_25(
        N_25_127));
    b8_1LbcQDr1_x_54_0 b9_1LbcgKeId (.mdiclink_reg({mdiclink_reg[322]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[54]}), .b4_nUAi({
        b4_nUAi[968], b4_nUAi[967], b4_nUAi[966]}), .b6_2ZTGIf({
        \b6_2ZTGIf[322] }));
    b8_1LbcQDr1_x_201_0 b9_1LbcgKGJp (.mdiclink_reg({mdiclink_reg[175]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[201]}), .b4_nUAi({
        b4_nUAi[526], b4_nUAi[525]}), .N_27(N_27_64), .N_25(N_25_64));
    b8_1LbcQDr1_x_17_0 b9_1LbcgKeUq (.mdiclink_reg({mdiclink_reg[359]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[17]}), .b4_nUAi({
        b4_nUAi[1079], b4_nUAi[1078], b4_nUAi[1077]}), .b6_2ZTGIf({
        \b6_2ZTGIf[359] }));
    b8_1LbcQDr1_x_351_0 b8_1LbcgKwU (.mdiclink_reg({mdiclink_reg[25]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[351]}), .b4_nUAi({
        b4_nUAi[77], b4_nUAi[76], b4_nUAi[75]}), .b6_2ZTGIf({
        \b6_2ZTGIf[25] }));
    b8_1LbcQDr1_x_311_0 b8_1LbcgKoU (.mdiclink_reg({mdiclink_reg[65]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[311]}), .b4_nUAi({
        b4_nUAi[197], b4_nUAi[196], b4_nUAi[195]}), .b6_2ZTGIf({
        \b6_2ZTGIf[65] }));
    b8_1LbcQDr1_x_163_0 b9_1LbcgKwSV (.mdiclink_reg({mdiclink_reg[213]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[163]}), .b4_nUAi({
        b4_nUAi[640], b4_nUAi[639]}), .N_27(N_27_77), .N_25(N_25_77));
    b8_1LbcQDr1_x_342_0 b8_1LbcgKeQ0 (.mdiclink_reg({mdiclink_reg[34]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[342]}), .b4_nUAi({
        b4_nUAi[104], b4_nUAi[103], b4_nUAi[102]}), .b6_2ZTGIf({
        \b6_2ZTGIf[34] }));
    b8_1LbcQDr1_x_212_0 b9_1LbcgKGAl (.mdiclink_reg({mdiclink_reg[164]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[212]}), .b4_nUAi({
        b4_nUAi[494], b4_nUAi[493], b4_nUAi[492]}), .b6_2ZTGIf({
        \b6_2ZTGIf[164] }));
    b8_1LbcQDr1_x_42_0 b9_1LbcgKeql (.mdiclink_reg({mdiclink_reg[334]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[42]}), .b4_nUAi({
        b4_nUAi[1003], b4_nUAi[1002]}), .N_27(N_27_123), .N_25(
        N_25_123));
    b8_1LbcQDr1_x_173_0 b9_1LbcgKwRV (.mdiclink_reg({mdiclink_reg[203]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[173]}), .b4_nUAi({
        b4_nUAi[610], b4_nUAi[609]}), .N_27(N_27_72), .N_25(N_25_72));
    b8_1LbcQDr1_x_210_0 b9_1LbcgKGA5 (.mdiclink_reg({mdiclink_reg[166]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[210]}), .b4_nUAi({
        b4_nUAi[500], b4_nUAi[499], b4_nUAi[498]}), .b6_2ZTGIf({
        \b6_2ZTGIf[166] }));
    b8_1LbcQDr1_x_312_0 b8_1LbcgKoQ0 (.mdiclink_reg({mdiclink_reg[64]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[312]}), .b4_nUAi({
        b4_nUAi[194], b4_nUAi[193], b4_nUAi[192]}), .b6_2ZTGIf({
        \b6_2ZTGIf[64] }));
    b8_1LbcQDr1_x_82_0 b9_1LbcgKwVl (.mdiclink_reg({mdiclink_reg[294]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[82]}), .b4_nUAi({
        b4_nUAi[884], b4_nUAi[883], b4_nUAi[882]}), .b6_2ZTGIf({
        \b6_2ZTGIf[294] }));
    b8_1LbcQDr1_x_146_0 b9_1LbcgKwqm (.mdiclink_reg({mdiclink_reg[230]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[146]}), .b4_nUAi({
        b4_nUAi[692], b4_nUAi[691], b4_nUAi[690]}), .b6_2ZTGIf({
        \b6_2ZTGIf[230] }));
    b8_1LbcQDr1_x_197_0 b9_1LbcgKGJq (.mdiclink_reg({mdiclink_reg[179]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[197]}), .b4_nUAi({
        b4_nUAi[539], b4_nUAi[538], b4_nUAi[537]}), .b6_2ZTGIf({
        \b6_2ZTGIf[179] }));
    b8_1LbcQDr1_x_125_0 b9_1LbcgKwUn (.mdiclink_reg({mdiclink_reg[251]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[125]}), .b4_nUAi({
        b4_nUAi[754], b4_nUAi[753]}), .N_27(N_27_90), .N_25(N_25_90));
    b8_1LbcQDr1_x_232_0 b9_1LbcgKGQl0 (.mdiclink_reg({
        mdiclink_reg[144]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[232]}), 
        .b4_nUAi({b4_nUAi[434], b4_nUAi[433], b4_nUAi[432]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[144] }));
    b8_1LbcQDr1_x_46_0 b9_1LbcgKeqm (.mdiclink_reg({mdiclink_reg[330]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[46]}), .b4_nUAi({
        b4_nUAi[992], b4_nUAi[991], b4_nUAi[990]}), .b6_2ZTGIf({
        \b6_2ZTGIf[330] }));
    b8_1LbcQDr1_x_107_0 b9_1LbcgKwAq (.mdiclink_reg({mdiclink_reg[269]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[107]}), .b4_nUAi({
        b4_nUAi[808], b4_nUAi[807]}), .N_27(N_27_98), .N_25(N_25_98));
    b8_1LbcQDr1_x_230_0 b9_1LbcgKGQ50 (.mdiclink_reg({
        mdiclink_reg[146]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[230]}), 
        .b4_nUAi({b4_nUAi[440], b4_nUAi[439], b4_nUAi[438]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[146] }));
    b8_1LbcQDr1_x_198_0 b9_1LbcgKGJS (.mdiclink_reg({mdiclink_reg[178]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[198]}), .b4_nUAi({
        b4_nUAi[536], b4_nUAi[535], b4_nUAi[534]}), .b6_2ZTGIf({
        \b6_2ZTGIf[178] }));
    b8_1LbcQDr1_x_109_0 b9_1LbcgKwAe (.mdiclink_reg({mdiclink_reg[267]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[109]}), .b4_nUAi({
        b4_nUAi[802], b4_nUAi[801]}), .N_27(N_27_96), .N_25(N_25_96));
    b8_1LbcQDr1_x_223_0 b9_1LbcgKGUV (.mdiclink_reg({mdiclink_reg[153]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[223]}), .b4_nUAi({
        b4_nUAi[461], b4_nUAi[460], b4_nUAi[459]}), .b6_2ZTGIf({
        \b6_2ZTGIf[153] }));
    b8_1LbcQDr1_x_199_0 b9_1LbcgKGJe (.mdiclink_reg({mdiclink_reg[177]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[199]}), .b4_nUAi({
        b4_nUAi[533], b4_nUAi[532], b4_nUAi[531]}), .b6_2ZTGIf({
        \b6_2ZTGIf[177] }));
    b8_1LbcQDr1_x_352_0 b8_1LbcgKwQ0 (.mdiclink_reg({mdiclink_reg[24]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[352]}), .b4_nUAi({
        b4_nUAi[74], b4_nUAi[73], b4_nUAi[72]}), .b6_2ZTGIf({
        \b6_2ZTGIf[24] }));
    b8_1LbcQDr1_x_127_0 b9_1LbcgKwQq0 (.mdiclink_reg({
        mdiclink_reg[249]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[127]}), 
        .b4_nUAi({b4_nUAi[749], b4_nUAi[748], b4_nUAi[747]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[249] }));
    b8_1LbcQDr1_x_158_0 b9_1LbcgKwSS (.mdiclink_reg({mdiclink_reg[218]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[158]}), .b4_nUAi({
        b4_nUAi[656], b4_nUAi[655], b4_nUAi[654]}), .b6_2ZTGIf({
        \b6_2ZTGIf[218] }));
    b8_1LbcQDr1_x_47_0 b9_1LbcgKeIq (.mdiclink_reg({mdiclink_reg[329]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[47]}), .b4_nUAi({
        b4_nUAi[989], b4_nUAi[988], b4_nUAi[987]}), .b6_2ZTGIf({
        \b6_2ZTGIf[329] }));
    b8_1LbcQDr1_x_354_0 b8_1LbcgKwI (.mdiclink_reg({mdiclink_reg[22]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[354]}), .b4_nUAi({
        b4_nUAi[68], b4_nUAi[67], b4_nUAi[66]}), .b6_2ZTGIf({
        \b6_2ZTGIf[22] }));
    b8_1LbcQDr1_x_314_0 b8_1LbcgKoI (.mdiclink_reg({mdiclink_reg[62]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[314]}), .b4_nUAi({
        b4_nUAi[187], b4_nUAi[186]}), .N_27(N_27_21), .N_25(N_25_21));
    b8_1LbcQDr1_x_168_0 b9_1LbcgKwRS (.mdiclink_reg({mdiclink_reg[208]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[168]}), .b4_nUAi({
        b4_nUAi[626], b4_nUAi[625], b4_nUAi[624]}), .b6_2ZTGIf({
        \b6_2ZTGIf[208] }));
    b8_1LbcQDr1_x_129_0 b9_1LbcgKwQe0 (.mdiclink_reg({
        mdiclink_reg[247]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[129]}), 
        .b4_nUAi({b4_nUAi[743], b4_nUAi[742], b4_nUAi[741]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[247] }));
    b8_1LbcQDr1_x_206_0 b9_1LbcgKGJm (.mdiclink_reg({mdiclink_reg[170]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[206]}), .b4_nUAi({
        b4_nUAi[512], b4_nUAi[511], b4_nUAi[510]}), .b6_2ZTGIf({
        \b6_2ZTGIf[170] }));
    b8_1LbcQDr1_x_94_0 b9_1LbcgKwnd (.mdiclink_reg({mdiclink_reg[282]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[94]}), .b4_nUAi({
        b4_nUAi[848], b4_nUAi[847], b4_nUAi[846]}), .b6_2ZTGIf({
        \b6_2ZTGIf[282] }));
    b8_1LbcQDr1_x_1_0 b9_1LbcgKeJp (.mdiclink_reg({mdiclink_reg[375]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[1]}), .b4_nUAi({
        b4_nUAi[1127], b4_nUAi[1126], b4_nUAi[1125]}), .b6_2ZTGIf({
        \b6_2ZTGIf[375] }));
    b8_1LbcQDr1_x_335_0 b8_1LbcgKES0 (.mdiclink_reg({mdiclink_reg[41]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[335]}), .b4_nUAi({
        b4_nUAi[125], b4_nUAi[124], b4_nUAi[123]}), .b6_2ZTGIf({
        \b6_2ZTGIf[41] }));
    b8_1LbcQDr1_x_298_0 b8_1LbcgKxn (.mdiclink_reg({mdiclink_reg[78]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[298]}), .b4_nUAi({
        b4_nUAi[235], b4_nUAi[234]}), .N_27(N_27_27), .N_25(N_25_27));
    b8_1LbcQDr1_x_358_0 b8_1LbcgKGn (.mdiclink_reg({mdiclink_reg[18]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[358]}), .b4_nUAi({
        b4_nUAi[56], b4_nUAi[55], b4_nUAi[54]}), .b6_2ZTGIf({
        \b6_2ZTGIf[18] }));
    b8_1LbcQDr1_x_155_0 b9_1LbcgKwIn (.mdiclink_reg({mdiclink_reg[221]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[155]}), .b4_nUAi({
        b4_nUAi[664], b4_nUAi[663]}), .N_27(N_27_80), .N_25(N_25_80));
    b8_1LbcQDr1_x_62_0 b9_1LbcgKeSl (.mdiclink_reg({mdiclink_reg[314]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[62]}), .b4_nUAi({
        b4_nUAi[944], b4_nUAi[943], b4_nUAi[942]}), .b6_2ZTGIf({
        \b6_2ZTGIf[314] }));
    b8_1LbcQDr1_x_38_0 b9_1LbcgKeqS (.mdiclink_reg({mdiclink_reg[338]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[38]}), .b4_nUAi({
        b4_nUAi[1016], b4_nUAi[1015], b4_nUAi[1014]}), .b6_2ZTGIf({
        \b6_2ZTGIf[338] }));
    b8_1LbcQDr1_x_289_0 b8_1LbcgKbJ (.mdiclink_reg({mdiclink_reg[87]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[289]}), .b4_nUAi({
        b4_nUAi[263], b4_nUAi[262], b4_nUAi[261]}), .b6_2ZTGIf({
        \b6_2ZTGIf[87] }));
    b8_1LbcQDr1_x_336_0 b8_1LbcgKER0 (.mdiclink_reg({mdiclink_reg[40]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[336]}), .b4_nUAi({
        b4_nUAi[122], b4_nUAi[121], b4_nUAi[120]}), .b6_2ZTGIf({
        \b6_2ZTGIf[40] }));
    b8_1LbcQDr1_x_340_0 b8_1LbcgKeA (.mdiclink_reg({mdiclink_reg[36]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[340]}), .b4_nUAi({
        b4_nUAi[110], b4_nUAi[109], b4_nUAi[108]}), .b6_2ZTGIf({
        \b6_2ZTGIf[36] }));
    b8_1LbcQDr1_x_166_0 b9_1LbcgKwSm (.mdiclink_reg({mdiclink_reg[210]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[166]}), .b4_nUAi({
        b4_nUAi[632], b4_nUAi[631], b4_nUAi[630]}), .b6_2ZTGIf({
        \b6_2ZTGIf[210] }));
    b8_1LbcQDr1_x_72_0 b9_1LbcgKeRl (.mdiclink_reg({mdiclink_reg[304]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[72]}), .b4_nUAi({
        b4_nUAi[914], b4_nUAi[913], b4_nUAi[912]}), .b6_2ZTGIf({
        \b6_2ZTGIf[304] }));
    b8_1LbcQDr1_x_318_0 b8_1LbcgKIn (.mdiclink_reg({mdiclink_reg[58]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[318]}), .b4_nUAi({
        b4_nUAi[176], b4_nUAi[175], b4_nUAi[174]}), .b6_2ZTGIf({
        \b6_2ZTGIf[58] }));
    b8_1LbcQDr1_x_176_0 b9_1LbcgKwRm (.mdiclink_reg({mdiclink_reg[200]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[176]}), .b4_nUAi({
        b4_nUAi[602], b4_nUAi[601], b4_nUAi[600]}), .b6_2ZTGIf({
        \b6_2ZTGIf[200] }));
    b8_1LbcQDr1_x_205_0 b9_1LbcgKGJn (.mdiclink_reg({mdiclink_reg[171]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[205]}), .b4_nUAi({
        b4_nUAi[514], b4_nUAi[513]}), .N_27(N_27_60), .N_25(N_25_60));
    b8_1LbcQDr1_x_253_0 b9_1LbcgKGIV (.mdiclink_reg({mdiclink_reg[123]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[253]}), .b4_nUAi({
        b4_nUAi[370], b4_nUAi[369]}), .N_27(N_27_42), .N_25(N_25_42));
    b8_1LbcQDr1_x_66_0 b9_1LbcgKeSm (.mdiclink_reg({mdiclink_reg[310]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[66]}), .b4_nUAi({
        b4_nUAi[932], b4_nUAi[931], b4_nUAi[930]}), .b6_2ZTGIf({
        \b6_2ZTGIf[310] }));
    b8_1LbcQDr1_x_84_0 b9_1LbcgKwVd (.mdiclink_reg({mdiclink_reg[292]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[84]}), .b4_nUAi({
        b4_nUAi[878], b4_nUAi[877], b4_nUAi[876]}), .b6_2ZTGIf({
        \b6_2ZTGIf[292] }));
    GND GND (.Y(GND_net_1));
    b8_1LbcQDr1_x_76_0 b9_1LbcgKeRm (.mdiclink_reg({mdiclink_reg[300]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[76]}), .b4_nUAi({
        b4_nUAi[901], b4_nUAi[900]}), .N_27(N_27_109), .N_25(N_25_109));
    b8_1LbcQDr1_x_297_0 b8_1LbcgKxV (.mdiclink_reg({mdiclink_reg[79]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[297]}), .b4_nUAi({
        b4_nUAi[238], b4_nUAi[237]}), .N_27(N_27_28), .N_25(N_25_28));
    b8_1LbcQDr1_x_357_0 b8_1LbcgKGV (.mdiclink_reg({mdiclink_reg[19]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[357]}), .b4_nUAi({
        b4_nUAi[59], b4_nUAi[58], b4_nUAi[57]}), .b6_2ZTGIf({
        \b6_2ZTGIf[19] }));
    b8_1LbcQDr1_x_4_0 b9_1LbcgKeJd (.mdiclink_reg({mdiclink_reg[372]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[4]}), .b4_nUAi({
        b4_nUAi[1117], b4_nUAi[1116]}), .N_27(N_27_139), .N_25(
        N_25_139));
    b8_1LbcQDr1_x_110_0 b9_1LbcgKwA5 (.mdiclink_reg({mdiclink_reg[266]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[110]}), .b4_nUAi({
        b4_nUAi[800], b4_nUAi[799], b4_nUAi[798]}), .b6_2ZTGIf({
        \b6_2ZTGIf[266] }));
    b8_1LbcQDr1_x_242_0 b9_1LbcgKGql (.mdiclink_reg({mdiclink_reg[134]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[242]}), .b4_nUAi({
        b4_nUAi[404], b4_nUAi[403], b4_nUAi[402]}), .b6_2ZTGIf({
        \b6_2ZTGIf[134] }));
    b8_1LbcQDr1_x_317_0 b8_1LbcgKIV (.mdiclink_reg({mdiclink_reg[59]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[317]}), .b4_nUAi({
        b4_nUAi[178], b4_nUAi[177]}), .N_27(N_27_18), .N_25(N_25_18));
    b8_1LbcQDr1_x_372_0 b7_1LbcgKE0 (.mdiclink_reg({mdiclink_reg[4]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[372]}), .b4_nUAi({
        b4_nUAi[14], b4_nUAi[13], b4_nUAi[12]}), .b6_2ZTGIf({
        \b6_2ZTGIf[4] }));
    b8_1LbcQDr1_x_240_0 b9_1LbcgKGq5 (.mdiclink_reg({mdiclink_reg[136]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[240]}), .b4_nUAi({
        b4_nUAi[410], b4_nUAi[409], b4_nUAi[408]}), .b6_2ZTGIf({
        \b6_2ZTGIf[136] }));
    b8_1LbcQDr1_x_122_0 b9_1LbcgKwUl (.mdiclink_reg({mdiclink_reg[254]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[122]}), .b4_nUAi({
        b4_nUAi[763], b4_nUAi[762]}), .N_27(N_27_93), .N_25(N_25_93));
    b8_1LbcQDr1_x_130_0 b9_1LbcgKwQ50 (.mdiclink_reg({
        mdiclink_reg[246]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[130]}), 
        .b4_nUAi({b4_nUAi[740], b4_nUAi[739], b4_nUAi[738]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[246] }));
    b8_1LbcQDr1_x_137_0 b9_1LbcgKwqq (.mdiclink_reg({mdiclink_reg[239]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[137]}), .b4_nUAi({
        b4_nUAi[718], b4_nUAi[717]}), .N_27(N_27_88), .N_25(N_25_88));
    b8_1LbcQDr1_x_93_0 b9_1LbcgKwnV (.mdiclink_reg({mdiclink_reg[283]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[93]}), .b4_nUAi({
        b4_nUAi[850], b4_nUAi[849]}), .N_27(N_27_102), .N_25(N_25_102));
    b8_1LbcQDr1_x_20_0 b9_1LbcgKeU5 (.mdiclink_reg({mdiclink_reg[356]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[20]}), .b4_nUAi({
        b4_nUAi[1070], b4_nUAi[1069], b4_nUAi[1068]}), .b6_2ZTGIf({
        \b6_2ZTGIf[356] }));
    b8_1LbcQDr1_x_139_0 b9_1LbcgKwqe (.mdiclink_reg({mdiclink_reg[237]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[139]}), .b4_nUAi({
        b4_nUAi[712], b4_nUAi[711]}), .N_27(N_27_86), .N_25(N_25_86));
    b8_1LbcQDr1_x_58_0 b9_1LbcgKeSS (.mdiclink_reg({mdiclink_reg[318]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[58]}), .b4_nUAi({
        b4_nUAi[955], b4_nUAi[954]}), .N_27(N_27_117), .N_25(N_25_117));
    b8_1LbcQDr1_x_68_0 b9_1LbcgKeRS (.mdiclink_reg({mdiclink_reg[308]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[68]}), .b4_nUAi({
        b4_nUAi[926], b4_nUAi[925], b4_nUAi[924]}), .b6_2ZTGIf({
        \b6_2ZTGIf[308] }));
    b8_1LbcQDr1_x_349_0 b8_1LbcgKwJ (.mdiclink_reg({mdiclink_reg[27]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[349]}), .b4_nUAi({
        b4_nUAi[82], b4_nUAi[81]}), .N_27(N_27_6), .N_25(N_25_6));
    b8_1LbcQDr1_x_83_0 b9_1LbcgKwVV (.mdiclink_reg({mdiclink_reg[293]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[83]}), .b4_nUAi({
        b4_nUAi[880], b4_nUAi[879]}), .N_27(N_27_107), .N_25(N_25_107));
    b8_1LbcQDr1_x_309_0 b8_1LbcgKoJ (.mdiclink_reg({mdiclink_reg[67]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[309]}), .b4_nUAi({
        b4_nUAi[203], b4_nUAi[202], b4_nUAi[201]}), .b6_2ZTGIf({
        \b6_2ZTGIf[67] }));
    b8_1LbcQDr1_x_152_0 b9_1LbcgKwIl (.mdiclink_reg({mdiclink_reg[224]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[152]}), .b4_nUAi({
        b4_nUAi[674], b4_nUAi[673], b4_nUAi[672]}), .b6_2ZTGIf({
        \b6_2ZTGIf[224] }));
    b8_1LbcQDr1_x_19_0 b9_1LbcgKeUe (.mdiclink_reg({mdiclink_reg[357]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[19]}), .b4_nUAi({
        b4_nUAi[1072], b4_nUAi[1071]}), .N_27(N_27_131), .N_25(
        N_25_131));
    b8_1LbcQDr1_x_262_0 b9_1LbcgKGSl (.mdiclink_reg({mdiclink_reg[114]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[262]}), .b4_nUAi({
        b4_nUAi[344], b4_nUAi[343], b4_nUAi[342]}), .b6_2ZTGIf({
        \b6_2ZTGIf[114] }));
    b8_1LbcQDr1_x_88_0 b9_1LbcgKwnS (.mdiclink_reg({mdiclink_reg[288]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[88]}), .b4_nUAi({
        b4_nUAi[866], b4_nUAi[865], b4_nUAi[864]}), .b6_2ZTGIf({
        \b6_2ZTGIf[288] }));
    b8_1LbcQDr1_x_280_0 b8_1LbcgKJA (.mdiclink_reg({mdiclink_reg[96]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[280]}), .b4_nUAi({
        b4_nUAi[290], b4_nUAi[289], b4_nUAi[288]}), .b6_2ZTGIf({
        \b6_2ZTGIf[96] }));
    b8_1LbcQDr1_x_260_0 b9_1LbcgKGS5 (.mdiclink_reg({mdiclink_reg[116]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[260]}), .b4_nUAi({
        b4_nUAi[350], b4_nUAi[349], b4_nUAi[348]}), .b6_2ZTGIf({
        \b6_2ZTGIf[116] }));
    b8_1LbcQDr1_x_105_0 b9_1LbcgKwJn (.mdiclink_reg({mdiclink_reg[271]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[105]}), .b4_nUAi({
        b4_nUAi[814], b4_nUAi[813]}), .N_27(N_27_100), .N_25(N_25_100));
    b8_1LbcQDr1_x_272_0 b9_1LbcgKGRl (.mdiclink_reg({mdiclink_reg[104]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[272]}), .b4_nUAi({
        b4_nUAi[314], b4_nUAi[313], b4_nUAi[312]}), .b6_2ZTGIf({
        \b6_2ZTGIf[104] }));
    b8_1LbcQDr1_x_343_0 b8_1LbcgKeq (.mdiclink_reg({mdiclink_reg[33]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[343]}), .b4_nUAi({
        b4_nUAi[101], b4_nUAi[100], b4_nUAi[99]}), .b6_2ZTGIf({
        \b6_2ZTGIf[33] }));
    b8_1LbcQDr1_x_270_0 b9_1LbcgKGR5 (.mdiclink_reg({mdiclink_reg[106]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[270]}), .b4_nUAi({
        b4_nUAi[320], b4_nUAi[319], b4_nUAi[318]}), .b6_2ZTGIf({
        \b6_2ZTGIf[106] }));
    b8_1LbcQDr1_x_50_0 b9_1LbcgKeI5 (.mdiclink_reg({mdiclink_reg[326]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[50]}), .b4_nUAi({
        b4_nUAi[980], b4_nUAi[979], b4_nUAi[978]}), .b6_2ZTGIf({
        \b6_2ZTGIf[326] }));
    b8_1LbcQDr1_x_124_0 b9_1LbcgKwUd (.mdiclink_reg({mdiclink_reg[252]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[124]}), .b4_nUAi({
        b4_nUAi[757], b4_nUAi[756]}), .N_27(N_27_91), .N_25(N_25_91));
    b8_1LbcQDr1_x_157_0 b9_1LbcgKwSq (.mdiclink_reg({mdiclink_reg[219]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[157]}), .b4_nUAi({
        b4_nUAi[658], b4_nUAi[657]}), .N_27(N_27_78), .N_25(N_25_78));
    b8_1LbcQDr1_x_203_0 b9_1LbcgKGJV (.mdiclink_reg({mdiclink_reg[173]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[203]}), .b4_nUAi({
        b4_nUAi[520], b4_nUAi[519]}), .N_27(N_27_62), .N_25(N_25_62));
    b8_1LbcQDr1_x_328_0 b8_1LbcgKEn0 (.mdiclink_reg({mdiclink_reg[48]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[328]}), .b4_nUAi({
        b4_nUAi[146], b4_nUAi[145], b4_nUAi[144]}), .b6_2ZTGIf({
        \b6_2ZTGIf[48] }));
    b8_1LbcQDr1_x_301_0 b8_1LbcgKxU (.mdiclink_reg({mdiclink_reg[75]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[301]}), .b4_nUAi({
        b4_nUAi[226], b4_nUAi[225]}), .N_27(N_27_24), .N_25(N_25_24));
    b8_1LbcQDr1_x_361_0 b8_1LbcgKGU (.mdiclink_reg({mdiclink_reg[15]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[361]}), .b4_nUAi({
        b4_nUAi[46], b4_nUAi[45]}), .N_27(N_27_4), .N_25(N_25_4));
    b8_1LbcQDr1_x_78_0 b9_1LbcgKwVS (.mdiclink_reg({mdiclink_reg[298]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[78]}), .b4_nUAi({
        b4_nUAi[896], b4_nUAi[895], b4_nUAi[894]}), .b6_2ZTGIf({
        \b6_2ZTGIf[298] }));
    b8_1LbcQDr1_x_167_0 b9_1LbcgKwRq (.mdiclink_reg({mdiclink_reg[209]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[167]}), .b4_nUAi({
        b4_nUAi[629], b4_nUAi[628], b4_nUAi[627]}), .b6_2ZTGIf({
        \b6_2ZTGIf[209] }));
    b8_1LbcQDr1_x_159_0 b9_1LbcgKwSe (.mdiclink_reg({mdiclink_reg[217]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[159]}), .b4_nUAi({
        b4_nUAi[653], b4_nUAi[652], b4_nUAi[651]}), .b6_2ZTGIf({
        \b6_2ZTGIf[217] }));
    b8_1LbcQDr1_x_369_0 b7_1LbcgKx (.mdiclink_reg({mdiclink_reg[7]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[369]}), .b4_nUAi({
        b4_nUAi[23], b4_nUAi[22], b4_nUAi[21]}), .b6_2ZTGIf({
        \b6_2ZTGIf[7] }));
    b8_1LbcQDr1_x_96_0 b9_1LbcgKwnm (.mdiclink_reg({mdiclink_reg[280]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[96]}), .b4_nUAi({
        b4_nUAi[842], b4_nUAi[841], b4_nUAi[840]}), .b6_2ZTGIf({
        \b6_2ZTGIf[280] }));
    b8_1LbcQDr1_x_140_0 b9_1LbcgKwq5 (.mdiclink_reg({mdiclink_reg[236]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[140]}), .b4_nUAi({
        b4_nUAi[709], b4_nUAi[708]}), .N_27(N_27_85), .N_25(N_25_85));
    b8_1LbcQDr1_x_13_0 b9_1LbcgKeAV (.mdiclink_reg({mdiclink_reg[363]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[13]}), .b4_nUAi({
        b4_nUAi[1090], b4_nUAi[1089]}), .N_27(N_27_132), .N_25(
        N_25_132));
    b8_1LbcQDr1_x_169_0 b9_1LbcgKwRe (.mdiclink_reg({mdiclink_reg[207]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[169]}), .b4_nUAi({
        b4_nUAi[622], b4_nUAi[621]}), .N_27(N_27_76), .N_25(N_25_76));
    b8_1LbcQDr1_x_321_0 b8_1LbcgKIU (.mdiclink_reg({mdiclink_reg[55]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[321]}), .b4_nUAi({
        b4_nUAi[167], b4_nUAi[166], b4_nUAi[165]}), .b6_2ZTGIf({
        \b6_2ZTGIf[55] }));
    b8_1LbcQDr1_x_49_0 b9_1LbcgKeIe (.mdiclink_reg({mdiclink_reg[327]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[49]}), .b4_nUAi({
        b4_nUAi[983], b4_nUAi[982], b4_nUAi[981]}), .b6_2ZTGIf({
        \b6_2ZTGIf[327] }));
    b8_1LbcQDr1_x_327_0 b8_1LbcgKEV0 (.mdiclink_reg({mdiclink_reg[49]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[327]}), .b4_nUAi({
        b4_nUAi[149], b4_nUAi[148], b4_nUAi[147]}), .b6_2ZTGIf({
        \b6_2ZTGIf[49] }));
    b8_1LbcQDr1_x_33_0 b9_1LbcgKeQV0 (.mdiclink_reg({mdiclink_reg[343]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[33]}), .b4_nUAi({
        b4_nUAi[1031], b4_nUAi[1030], b4_nUAi[1029]}), .b6_2ZTGIf({
        \b6_2ZTGIf[343] }));
    b8_1LbcQDr1_x_25_0 b9_1LbcgKeUn (.mdiclink_reg({mdiclink_reg[351]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[25]}), .b4_nUAi({
        b4_nUAi[1054], b4_nUAi[1053]}), .N_27(N_27_130), .N_25(
        N_25_130));
    VCC VCC (.Y(VCC_net_1));
    b8_1LbcQDr1_x_86_0 b9_1LbcgKwVm (.mdiclink_reg({mdiclink_reg[290]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[86]}), .b4_nUAi({
        b4_nUAi[872], b4_nUAi[871], b4_nUAi[870]}), .b6_2ZTGIf({
        \b6_2ZTGIf[290] }));
    b8_1LbcQDr1_x_332_0 b8_1LbcgKEQ0 (.mdiclink_reg({mdiclink_reg[44]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[332]}), .b4_nUAi({
        b4_nUAi[133], b4_nUAi[132]}), .N_27(N_27_13), .N_25(N_25_13));
    b8_1LbcQDr1_x_154_0 b9_1LbcgKwId (.mdiclink_reg({mdiclink_reg[222]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[154]}), .b4_nUAi({
        b4_nUAi[667], b4_nUAi[666]}), .N_27(N_27_81), .N_25(N_25_81));
    b8_1LbcQDr1_x_345_0 b8_1LbcgKeS (.mdiclink_reg({mdiclink_reg[31]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[345]}), .b4_nUAi({
        b4_nUAi[94], b4_nUAi[93]}), .N_27(N_27_10), .N_25(N_25_10));
    b8_1LbcQDr1_x_111_0 b9_1LbcgKwAp (.mdiclink_reg({mdiclink_reg[265]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[111]}), .b4_nUAi({
        b4_nUAi[797], b4_nUAi[796], b4_nUAi[795]}), .b6_2ZTGIf({
        \b6_2ZTGIf[265] }));
    b8_1LbcQDr1_x_304_0 b8_1LbcgKxI (.mdiclink_reg({mdiclink_reg[72]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[304]}), .b4_nUAi({
        b4_nUAi[218], b4_nUAi[217], b4_nUAi[216]}), .b6_2ZTGIf({
        \b6_2ZTGIf[72] }));
    b8_1LbcQDr1_x_364_0 b8_1LbcgKGI (.mdiclink_reg({mdiclink_reg[12]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[364]}), .b4_nUAi({
        b4_nUAi[37], b4_nUAi[36]}), .N_27(N_27_1), .N_25(N_25_1));
    b8_1LbcQDr1_x_346_0 b8_1LbcgKeR (.mdiclink_reg({mdiclink_reg[30]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[346]}), .b4_nUAi({
        b4_nUAi[91], b4_nUAi[90]}), .N_27(N_27_9), .N_25(N_25_9));
    b8_1LbcQDr1_x_214_0 b9_1LbcgKGAd (.mdiclink_reg({mdiclink_reg[162]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[214]}), .b4_nUAi({
        b4_nUAi[488], b4_nUAi[487], b4_nUAi[486]}), .b6_2ZTGIf({
        \b6_2ZTGIf[162] }));
    b8_1LbcQDr1_x_123_0 b9_1LbcgKwUV (.mdiclink_reg({mdiclink_reg[253]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[123]}), .b4_nUAi({
        b4_nUAi[760], b4_nUAi[759]}), .N_27(N_27_92), .N_25(N_25_92));
    b8_1LbcQDr1_x_324_0 b8_1LbcgKII (.mdiclink_reg({mdiclink_reg[52]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[324]}), .b4_nUAi({
        b4_nUAi[158], b4_nUAi[157], b4_nUAi[156]}), .b6_2ZTGIf({
        \b6_2ZTGIf[52] }));
    b8_1LbcQDr1_x_131_0 b9_1LbcgKwQp0 (.mdiclink_reg({
        mdiclink_reg[245]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[131]}), 
        .b4_nUAi({b4_nUAi[736], b4_nUAi[735]}), .N_27(N_27_89), .N_25(
        N_25_89));
    b8_1LbcQDr1_x_102_0 b9_1LbcgKwJl (.mdiclink_reg({mdiclink_reg[274]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[102]}), .b4_nUAi({
        b4_nUAi[824], b4_nUAi[823], b4_nUAi[822]}), .b6_2ZTGIf({
        \b6_2ZTGIf[274] }));
    b8_1LbcQDr1_x_234_0 b9_1LbcgKGQd0 (.mdiclink_reg({
        mdiclink_reg[142]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[234]}), 
        .b4_nUAi({b4_nUAi[427], b4_nUAi[426]}), .N_27(N_27_51), .N_25(
        N_25_51));
    b8_1LbcQDr1_x_160_0 b9_1LbcgKwS5 (.mdiclink_reg({mdiclink_reg[216]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[160]}), .b4_nUAi({
        b4_nUAi[650], b4_nUAi[649], b4_nUAi[648]}), .b6_2ZTGIf({
        \b6_2ZTGIf[216] }));
    b8_1LbcQDr1_x_283_0 b8_1LbcgKJq (.mdiclink_reg({mdiclink_reg[93]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[283]}), .b4_nUAi({
        b4_nUAi[280], b4_nUAi[279]}), .N_27(N_27_32), .N_25(N_25_32));
    b8_1LbcQDr1_x_370_0 b7_1LbcgKo (.mdiclink_reg({mdiclink_reg[6]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[370]}), .b4_nUAi({
        b4_nUAi[20], b4_nUAi[19], b4_nUAi[18]}), .b6_2ZTGIf({
        \b6_2ZTGIf[6] }));
    b8_1LbcQDr1_x_170_0 b9_1LbcgKwR5 (.mdiclink_reg({mdiclink_reg[206]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[170]}), .b4_nUAi({
        b4_nUAi[619], b4_nUAi[618]}), .N_27(N_27_75), .N_25(N_25_75));
    b8_1LbcQDr1_x_55_0 b9_1LbcgKeIn (.mdiclink_reg({mdiclink_reg[321]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[55]}), .b4_nUAi({
        b4_nUAi[965], b4_nUAi[964], b4_nUAi[963]}), .b6_2ZTGIf({
        \b6_2ZTGIf[321] }));
    b8_1LbcQDr1_x_0_0 b9_1LbcgKeJ5 (.mdiclink_reg({mdiclink_reg[376]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[0]}), .b4_nUAi({
        b4_nUAi[1129], b4_nUAi[1128]}), .N_27(N_27_141), .N_25(
        N_25_141));
    b8_1LbcQDr1_x_211_0 b9_1LbcgKGAp (.mdiclink_reg({mdiclink_reg[165]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[211]}), .b4_nUAi({
        b4_nUAi[496], b4_nUAi[495]}), .N_27(N_27_59), .N_25(N_25_59));
    b8_1LbcQDr1_x_192_0 b9_1LbcgKGnl (.mdiclink_reg({mdiclink_reg[184]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[192]}), .b4_nUAi({
        b4_nUAi[554], b4_nUAi[553], b4_nUAi[552]}), .b6_2ZTGIf({
        \b6_2ZTGIf[184] }));
    b8_1LbcQDr1_x_118_0 b9_1LbcgKwUS (.mdiclink_reg({mdiclink_reg[258]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[118]}), .b4_nUAi({
        b4_nUAi[776], b4_nUAi[775], b4_nUAi[774]}), .b6_2ZTGIf({
        \b6_2ZTGIf[258] }));
    b8_1LbcQDr1_x_190_0 b9_1LbcgKGn5 (.mdiclink_reg({mdiclink_reg[186]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[190]}), .b4_nUAi({
        b4_nUAi[560], b4_nUAi[559], b4_nUAi[558]}), .b6_2ZTGIf({
        \b6_2ZTGIf[186] }));
    b8_1LbcQDr1_x_153_0 b9_1LbcgKwIV (.mdiclink_reg({mdiclink_reg[223]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[153]}), .b4_nUAi({
        b4_nUAi[670], b4_nUAi[669]}), .N_27(N_27_82), .N_25(N_25_82));
    b8_1LbcQDr1_x_43_0 b9_1LbcgKeqV (.mdiclink_reg({mdiclink_reg[333]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[43]}), .b4_nUAi({
        b4_nUAi[1000], b4_nUAi[999]}), .N_27(N_27_122), .N_25(N_25_122)
        );
    b8_1LbcQDr1_x_231_0 b9_1LbcgKGQp0 (.mdiclink_reg({
        mdiclink_reg[145]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[231]}), 
        .b4_nUAi({b4_nUAi[437], b4_nUAi[436], b4_nUAi[435]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[145] }));
    b8_1LbcQDr1_x_207_0 b9_1LbcgKGAq (.mdiclink_reg({mdiclink_reg[169]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[207]}), .b4_nUAi({
        b4_nUAi[509], b4_nUAi[508], b4_nUAi[507]}), .b6_2ZTGIf({
        \b6_2ZTGIf[169] }));
    b8_1LbcQDr1_x_87_0 b9_1LbcgKwnq (.mdiclink_reg({mdiclink_reg[289]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[87]}), .b4_nUAi({
        b4_nUAi[869], b4_nUAi[868], b4_nUAi[867]}), .b6_2ZTGIf({
        \b6_2ZTGIf[289] }));
    b8_1LbcQDr1_x_331_0 b8_1LbcgKEU0 (.mdiclink_reg({mdiclink_reg[45]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[331]}), .b4_nUAi({
        b4_nUAi[136], b4_nUAi[135]}), .N_27(N_27_14), .N_25(N_25_14));
    b8_1LbcQDr1_x_182_0 b9_1LbcgKGVl (.mdiclink_reg({mdiclink_reg[194]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[182]}), .b4_nUAi({
        b4_nUAi[584], b4_nUAi[583], b4_nUAi[582]}), .b6_2ZTGIf({
        \b6_2ZTGIf[194] }));
    b8_1LbcQDr1_x_208_0 b9_1LbcgKGAS (.mdiclink_reg({mdiclink_reg[168]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[208]}), .b4_nUAi({
        b4_nUAi[506], b4_nUAi[505], b4_nUAi[504]}), .b6_2ZTGIf({
        \b6_2ZTGIf[168] }));
    b8_1LbcQDr1_x_22_0 b9_1LbcgKeUl (.mdiclink_reg({mdiclink_reg[354]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[22]}), .b4_nUAi({
        b4_nUAi[1064], b4_nUAi[1063], b4_nUAi[1062]}), .b6_2ZTGIf({
        \b6_2ZTGIf[354] }));
    b8_1LbcQDr1_x_89_0 b9_1LbcgKwne (.mdiclink_reg({mdiclink_reg[287]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[89]}), .b4_nUAi({
        b4_nUAi[862], b4_nUAi[861]}), .N_27(N_27_106), .N_25(N_25_106));
    b8_1LbcQDr1_x_180_0 b9_1LbcgKGV5 (.mdiclink_reg({mdiclink_reg[196]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[180]}), .b4_nUAi({
        b4_nUAi[590], b4_nUAi[589], b4_nUAi[588]}), .b6_2ZTGIf({
        \b6_2ZTGIf[196] }));
    b8_1LbcQDr1_x_126_0 b9_1LbcgKwUm (.mdiclink_reg({mdiclink_reg[250]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[126]}), .b4_nUAi({
        b4_nUAi[752], b4_nUAi[751], b4_nUAi[750]}), .b6_2ZTGIf({
        \b6_2ZTGIf[250] }));
    b8_1LbcQDr1_x_227_0 b9_1LbcgKGQq0 (.mdiclink_reg({
        mdiclink_reg[149]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[227]}), 
        .b4_nUAi({b4_nUAi[448], b4_nUAi[447]}), .N_27(N_27_53), .N_25(
        N_25_53));
    b8_1LbcQDr1_x_209_0 b9_1LbcgKGAe (.mdiclink_reg({mdiclink_reg[167]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[209]}), .b4_nUAi({
        b4_nUAi[503], b4_nUAi[502], b4_nUAi[501]}), .b6_2ZTGIf({
        \b6_2ZTGIf[167] }));
    b8_1LbcQDr1_x_285_0 b8_1LbcgKJS (.mdiclink_reg({mdiclink_reg[91]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[285]}), .b4_nUAi({
        b4_nUAi[274], b4_nUAi[273]}), .N_27(N_27_30), .N_25(N_25_30));
    b8_1LbcQDr1_x_26_0 b9_1LbcgKeUm (.mdiclink_reg({mdiclink_reg[350]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[26]}), .b4_nUAi({
        b4_nUAi[1051], b4_nUAi[1050]}), .N_27(N_27_129), .N_25(
        N_25_129));
    b8_1LbcQDr1_x_371_0 b7_1LbcgKI (.mdiclink_reg({mdiclink_reg[5]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[371]}), .b4_nUAi({
        b4_nUAi[16], b4_nUAi[15]}), .N_27(N_27), .N_25(N_25));
    b8_1LbcQDr1_x_228_0 b9_1LbcgKGQS0 (.mdiclink_reg({
        mdiclink_reg[148]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[228]}), 
        .b4_nUAi({b4_nUAi[446], b4_nUAi[445], b4_nUAi[444]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[148] }));
    b8_1LbcQDr1_x_77_0 b9_1LbcgKwVq (.mdiclink_reg({mdiclink_reg[299]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[77]}), .b4_nUAi({
        b4_nUAi[898], b4_nUAi[897]}), .N_27(N_27_108), .N_25(N_25_108));
    b8_1LbcQDr1_x_286_0 b8_1LbcgKJR (.mdiclink_reg({mdiclink_reg[90]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[286]}), .b4_nUAi({
        b4_nUAi[272], b4_nUAi[271], b4_nUAi[270]}), .b6_2ZTGIf({
        \b6_2ZTGIf[90] }));
    b8_1LbcQDr1_x_141_0 b9_1LbcgKwqp (.mdiclink_reg({mdiclink_reg[235]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[141]}), .b4_nUAi({
        b4_nUAi[706], b4_nUAi[705]}), .N_27(N_27_84), .N_25(N_25_84));
    b8_1LbcQDr1_x_104_0 b9_1LbcgKwJd (.mdiclink_reg({mdiclink_reg[272]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[104]}), .b4_nUAi({
        b4_nUAi[818], b4_nUAi[817], b4_nUAi[816]}), .b6_2ZTGIf({
        \b6_2ZTGIf[272] }));
    b8_1LbcQDr1_x_216_0 b9_1LbcgKGAm (.mdiclink_reg({mdiclink_reg[160]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[216]}), .b4_nUAi({
        b4_nUAi[482], b4_nUAi[481], b4_nUAi[480]}), .b6_2ZTGIf({
        \b6_2ZTGIf[160] }));
    b8_1LbcQDr1_x_148_0 b9_1LbcgKwIS (.mdiclink_reg({mdiclink_reg[228]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[148]}), .b4_nUAi({
        b4_nUAi[686], b4_nUAi[685], b4_nUAi[684]}), .b6_2ZTGIf({
        \b6_2ZTGIf[228] }));
    b8_1LbcQDr1_x_244_0 b9_1LbcgKGqd (.mdiclink_reg({mdiclink_reg[132]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[244]}), .b4_nUAi({
        b4_nUAi[398], b4_nUAi[397], b4_nUAi[396]}), .b6_2ZTGIf({
        \b6_2ZTGIf[132] }));
    b8_1LbcQDr1_x_79_0 b9_1LbcgKwVe (.mdiclink_reg({mdiclink_reg[297]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[79]}), .b4_nUAi({
        b4_nUAi[893], b4_nUAi[892], b4_nUAi[891]}), .b6_2ZTGIf({
        \b6_2ZTGIf[297] }));
    b8_1LbcQDr1_x_229_0 b9_1LbcgKGQe0 (.mdiclink_reg({
        mdiclink_reg[147]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[229]}), 
        .b4_nUAi({b4_nUAi[443], b4_nUAi[442], b4_nUAi[441]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[147] }));
    b8_1LbcQDr1_x_299_0 b8_1LbcgKxJ (.mdiclink_reg({mdiclink_reg[77]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[299]}), .b4_nUAi({
        b4_nUAi[232], b4_nUAi[231]}), .N_27(N_27_26), .N_25(N_25_26));
    b8_1LbcQDr1_x_359_0 b8_1LbcgKGJ (.mdiclink_reg({mdiclink_reg[17]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[359]}), .b4_nUAi({
        b4_nUAi[53], b4_nUAi[52], b4_nUAi[51]}), .b6_2ZTGIf({
        \b6_2ZTGIf[17] }));
    b8_1LbcQDr1_x_322_0 b8_1LbcgKIQ0 (.mdiclink_reg({mdiclink_reg[54]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[322]}), .b4_nUAi({
        b4_nUAi[164], b4_nUAi[163], b4_nUAi[162]}), .b6_2ZTGIf({
        \b6_2ZTGIf[54] }));
    b8_1LbcQDr1_x_374_0 b7_1LbcgKw (.mdiclink_reg({mdiclink_reg[2]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[374]}), .b4_nUAi({b4_nUAi[8], 
        b4_nUAi[7], b4_nUAi[6]}), .b6_2ZTGIf({\b6_2ZTGIf[2] }));
    b8_1LbcQDr1_x_11_0 b9_1LbcgKeAp (.mdiclink_reg({mdiclink_reg[365]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[11]}), .b4_nUAi({
        b4_nUAi[1096], b4_nUAi[1095]}), .N_27(N_27_134), .N_25(
        N_25_134));
    b8_1LbcQDr1_x_319_0 b8_1LbcgKIJ (.mdiclink_reg({mdiclink_reg[57]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[319]}), .b4_nUAi({
        b4_nUAi[173], b4_nUAi[172], b4_nUAi[171]}), .b6_2ZTGIf({
        \b6_2ZTGIf[57] }));
    b8_1LbcQDr1_x_236_0 b9_1LbcgKGQm0 (.mdiclink_reg({
        mdiclink_reg[140]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[236]}), 
        .b4_nUAi({b4_nUAi[421], b4_nUAi[420]}), .N_27(N_27_49), .N_25(
        N_25_49));
    b8_1LbcQDr1_x_338_0 b8_1LbcgKen (.mdiclink_reg({mdiclink_reg[38]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[338]}), .b4_nUAi({
        b4_nUAi[116], b4_nUAi[115], b4_nUAi[114]}), .b6_2ZTGIf({
        \b6_2ZTGIf[38] }));
    b8_1LbcQDr1_x_290_0 b8_1LbcgKbA (.mdiclink_reg({mdiclink_reg[86]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[290]}), .b4_nUAi({
        b4_nUAi[260], b4_nUAi[259], b4_nUAi[258]}), .b6_2ZTGIf({
        \b6_2ZTGIf[86] }));
    b8_1LbcQDr1_x_63_0 b9_1LbcgKeSV (.mdiclink_reg({mdiclink_reg[313]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[63]}), .b4_nUAi({
        b4_nUAi[941], b4_nUAi[940], b4_nUAi[939]}), .b6_2ZTGIf({
        \b6_2ZTGIf[313] }));
    b8_1LbcQDr1_x_334_0 b8_1LbcgKEI0 (.mdiclink_reg({mdiclink_reg[42]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[334]}), .b4_nUAi({
        b4_nUAi[128], b4_nUAi[127], b4_nUAi[126]}), .b6_2ZTGIf({
        \b6_2ZTGIf[42] }));
    b8_1LbcQDr1_x_52_0 b9_1LbcgKeIl (.mdiclink_reg({mdiclink_reg[324]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[52]}), .b4_nUAi({
        b4_nUAi[974], b4_nUAi[973], b4_nUAi[972]}), .b6_2ZTGIf({
        \b6_2ZTGIf[324] }));
    b8_1LbcQDr1_x_73_0 b9_1LbcgKeRV (.mdiclink_reg({mdiclink_reg[303]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[73]}), .b4_nUAi({
        b4_nUAi[910], b4_nUAi[909]}), .N_27(N_27_112), .N_25(N_25_112));
    b8_1LbcQDr1_x_31_0 b9_1LbcgKeQp0 (.mdiclink_reg({mdiclink_reg[345]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[31]}), .b4_nUAi({
        b4_nUAi[1037], b4_nUAi[1036], b4_nUAi[1035]}), .b6_2ZTGIf({
        \b6_2ZTGIf[345] }));
    b8_1LbcQDr1_x_156_0 b9_1LbcgKwIm (.mdiclink_reg({mdiclink_reg[220]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[156]}), .b4_nUAi({
        b4_nUAi[661], b4_nUAi[660]}), .N_27(N_27_79), .N_25(N_25_79));
    b8_1LbcQDr1_x_215_0 b9_1LbcgKGAn (.mdiclink_reg({mdiclink_reg[161]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[215]}), .b4_nUAi({
        b4_nUAi[485], b4_nUAi[484], b4_nUAi[483]}), .b6_2ZTGIf({
        \b6_2ZTGIf[161] }));
    b8_1LbcQDr1_x_5_0 b9_1LbcgKeJn (.mdiclink_reg({mdiclink_reg[371]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[5]}), .b4_nUAi({
        b4_nUAi[1115], b4_nUAi[1114], b4_nUAi[1113]}), .b6_2ZTGIf({
        \b6_2ZTGIf[371] }));
    b8_1LbcQDr1_x_18_0 b9_1LbcgKeUS (.mdiclink_reg({mdiclink_reg[358]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[18]}), .b4_nUAi({
        b4_nUAi[1076], b4_nUAi[1075], b4_nUAi[1074]}), .b6_2ZTGIf({
        \b6_2ZTGIf[358] }));
    b8_1LbcQDr1_x_241_0 b9_1LbcgKGqp (.mdiclink_reg({mdiclink_reg[135]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[241]}), .b4_nUAi({
        b4_nUAi[407], b4_nUAi[406], b4_nUAi[405]}), .b6_2ZTGIf({
        \b6_2ZTGIf[135] }));
    b8_1LbcQDr1_x_56_0 b9_1LbcgKeIm (.mdiclink_reg({mdiclink_reg[320]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[56]}), .b4_nUAi({
        b4_nUAi[962], b4_nUAi[961], b4_nUAi[960]}), .b6_2ZTGIf({
        \b6_2ZTGIf[320] }));
    b8_1LbcQDr1_x_14_0 b9_1LbcgKeAd (.mdiclink_reg({mdiclink_reg[362]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[14]}), .b4_nUAi({
        b4_nUAi[1088], b4_nUAi[1087], b4_nUAi[1086]}), .b6_2ZTGIf({
        \b6_2ZTGIf[362] }));
    b8_1LbcQDr1_x_337_0 b8_1LbcgKeV (.mdiclink_reg({mdiclink_reg[39]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[337]}), .b4_nUAi({
        b4_nUAi[119], b4_nUAi[118], b4_nUAi[117]}), .b6_2ZTGIf({
        \b6_2ZTGIf[39] }));
    b8_1LbcQDr1_x_90_0 b9_1LbcgKwn5 (.mdiclink_reg({mdiclink_reg[286]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[90]}), .b4_nUAi({
        b4_nUAi[859], b4_nUAi[858]}), .N_27(N_27_105), .N_25(N_25_105));
    b8_1LbcQDr1_x_235_0 b9_1LbcgKGQn0 (.mdiclink_reg({
        mdiclink_reg[141]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[235]}), 
        .b4_nUAi({b4_nUAi[424], b4_nUAi[423]}), .N_27(N_27_50), .N_25(
        N_25_50));
    b8_1LbcQDr1_x_161_0 b9_1LbcgKwSp (.mdiclink_reg({mdiclink_reg[215]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[161]}), .b4_nUAi({
        b4_nUAi[647], b4_nUAi[646], b4_nUAi[645]}), .b6_2ZTGIf({
        \b6_2ZTGIf[215] }));
    b8_1LbcQDr1_x_103_0 b9_1LbcgKwJV (.mdiclink_reg({mdiclink_reg[273]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[103]}), .b4_nUAi({
        b4_nUAi[821], b4_nUAi[820], b4_nUAi[819]}), .b6_2ZTGIf({
        \b6_2ZTGIf[273] }));
    b8_1LbcQDr1_x_34_0 b9_1LbcgKeQd0 (.mdiclink_reg({mdiclink_reg[342]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[34]}), .b4_nUAi({
        b4_nUAi[1028], b4_nUAi[1027], b4_nUAi[1026]}), .b6_2ZTGIf({
        \b6_2ZTGIf[342] }));
    b8_1LbcQDr1_x_237_0 b9_1LbcgKGqq (.mdiclink_reg({mdiclink_reg[139]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[237]}), .b4_nUAi({
        b4_nUAi[418], b4_nUAi[417]}), .N_27(N_27_48), .N_25(N_25_48));
    b8_1LbcQDr1_x_264_0 b9_1LbcgKGSd (.mdiclink_reg({mdiclink_reg[112]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[264]}), .b4_nUAi({
        b4_nUAi[338], b4_nUAi[337], b4_nUAi[336]}), .b6_2ZTGIf({
        \b6_2ZTGIf[112] }));
    b8_1LbcQDr1_x_171_0 b9_1LbcgKwRp (.mdiclink_reg({mdiclink_reg[205]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[171]}), .b4_nUAi({
        b4_nUAi[616], b4_nUAi[615]}), .N_27(N_27_74), .N_25(N_25_74));
    b8_1LbcQDr1_x_80_0 b9_1LbcgKwV5 (.mdiclink_reg({mdiclink_reg[296]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[80]}), .b4_nUAi({
        b4_nUAi[890], b4_nUAi[889], b4_nUAi[888]}), .b6_2ZTGIf({
        \b6_2ZTGIf[296] }));
    b8_1LbcQDr1_x_222_0 b9_1LbcgKGUl (.mdiclink_reg({mdiclink_reg[154]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[222]}), .b4_nUAi({
        b4_nUAi[464], b4_nUAi[463], b4_nUAi[462]}), .b6_2ZTGIf({
        \b6_2ZTGIf[154] }));
    b8_1LbcQDr1_x_274_0 b9_1LbcgKGRd (.mdiclink_reg({mdiclink_reg[102]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[274]}), .b4_nUAi({
        b4_nUAi[308], b4_nUAi[307], b4_nUAi[306]}), .b6_2ZTGIf({
        \b6_2ZTGIf[102] }));
    b8_1LbcQDr1_x_238_0 b9_1LbcgKGqS (.mdiclink_reg({mdiclink_reg[138]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[238]}), .b4_nUAi({
        b4_nUAi[416], b4_nUAi[415], b4_nUAi[414]}), .b6_2ZTGIf({
        \b6_2ZTGIf[138] }));
    b8_1LbcQDr1_x_220_0 b9_1LbcgKGU5 (.mdiclink_reg({mdiclink_reg[156]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[220]}), .b4_nUAi({
        b4_nUAi[469], b4_nUAi[468]}), .N_27(N_27_55), .N_25(N_25_55));
    b8_1LbcQDr1_x_239_0 b9_1LbcgKGqe (.mdiclink_reg({mdiclink_reg[137]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[239]}), .b4_nUAi({
        b4_nUAi[413], b4_nUAi[412], b4_nUAi[411]}), .b6_2ZTGIf({
        \b6_2ZTGIf[137] }));
    b8_1LbcQDr1_x_48_0 b9_1LbcgKeIS (.mdiclink_reg({mdiclink_reg[328]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[48]}), .b4_nUAi({
        b4_nUAi[986], b4_nUAi[985], b4_nUAi[984]}), .b6_2ZTGIf({
        \b6_2ZTGIf[328] }));
    b8_1LbcQDr1_x_117_0 b9_1LbcgKwUq (.mdiclink_reg({mdiclink_reg[259]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[117]}), .b4_nUAi({
        b4_nUAi[779], b4_nUAi[778], b4_nUAi[777]}), .b6_2ZTGIf({
        \b6_2ZTGIf[259] }));
    b8_1LbcQDr1_x_7_0 b9_1LbcgKeAq (.mdiclink_reg({mdiclink_reg[369]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[7]}), .b4_nUAi({
        b4_nUAi[1109], b4_nUAi[1108], b4_nUAi[1107]}), .b6_2ZTGIf({
        \b6_2ZTGIf[369] }));
    b8_1LbcQDr1_x_350_0 b8_1LbcgKwA (.mdiclink_reg({mdiclink_reg[26]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[350]}), .b4_nUAi({
        b4_nUAi[80], b4_nUAi[79], b4_nUAi[78]}), .b6_2ZTGIf({
        \b6_2ZTGIf[26] }));
    b8_1LbcQDr1_x_376_0 b7_1LbcgKF (.mdiclink_reg({mdiclink_reg[0]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[376]}), .b4_nUAi({b4_nUAi[2], 
        b4_nUAi[1], b4_nUAi[0]}), .b6_2ZTGIf({\b6_2ZTGIf[0] }));
    b8_1LbcQDr1_x_246_0 b9_1LbcgKGqm (.mdiclink_reg({mdiclink_reg[130]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[246]}), .b4_nUAi({
        b4_nUAi[392], b4_nUAi[391], b4_nUAi[390]}), .b6_2ZTGIf({
        \b6_2ZTGIf[130] }));
    b8_1LbcQDr1_x_310_0 b8_1LbcgKoA (.mdiclink_reg({mdiclink_reg[66]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[310]}), .b4_nUAi({
        b4_nUAi[200], b4_nUAi[199], b4_nUAi[198]}), .b6_2ZTGIf({
        \b6_2ZTGIf[66] }));
    b8_1LbcQDr1_x_119_0 b9_1LbcgKwUe (.mdiclink_reg({mdiclink_reg[257]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[119]}), .b4_nUAi({
        b4_nUAi[773], b4_nUAi[772], b4_nUAi[771]}), .b6_2ZTGIf({
        \b6_2ZTGIf[257] }));
    b8_1LbcQDr1_x_98_0 b9_1LbcgKwJS (.mdiclink_reg({mdiclink_reg[278]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[98]}), .b4_nUAi({
        b4_nUAi[836], b4_nUAi[835], b4_nUAi[834]}), .b6_2ZTGIf({
        \b6_2ZTGIf[278] }));
    b8_1LbcQDr1_x_261_0 b9_1LbcgKGSp (.mdiclink_reg({mdiclink_reg[115]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[261]}), .b4_nUAi({
        b4_nUAi[347], b4_nUAi[346], b4_nUAi[345]}), .b6_2ZTGIf({
        \b6_2ZTGIf[115] }));
    b8_1LbcQDr1_x_271_0 b9_1LbcgKGRp (.mdiclink_reg({mdiclink_reg[105]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[271]}), .b4_nUAi({
        b4_nUAi[317], b4_nUAi[316], b4_nUAi[315]}), .b6_2ZTGIf({
        \b6_2ZTGIf[105] }));
    b8_1LbcQDr1_x_41_0 b9_1LbcgKeqp (.mdiclink_reg({mdiclink_reg[335]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[41]}), .b4_nUAi({
        b4_nUAi[1006], b4_nUAi[1005]}), .N_27(N_27_124), .N_25(
        N_25_124));
    b8_1LbcQDr1_x_278_0 b8_1LbcgKJn (.mdiclink_reg({mdiclink_reg[98]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[278]}), .b4_nUAi({
        b4_nUAi[296], b4_nUAi[295], b4_nUAi[294]}), .b6_2ZTGIf({
        \b6_2ZTGIf[98] }));
    b8_1LbcQDr1_x_27_0 b9_1LbcgKeQq0 (.mdiclink_reg({mdiclink_reg[349]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[27]}), .b4_nUAi({
        b4_nUAi[1048], b4_nUAi[1047]}), .N_27(N_27_128), .N_25(
        N_25_128));
    b8_1LbcQDr1_x_293_0 b8_1LbcgKbq (.mdiclink_reg({mdiclink_reg[83]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[293]}), .b4_nUAi({
        b4_nUAi[251], b4_nUAi[250], b4_nUAi[249]}), .b6_2ZTGIf({
        \b6_2ZTGIf[83] }));
    b8_1LbcQDr1_x_115_0 b9_1LbcgKwAn (.mdiclink_reg({mdiclink_reg[261]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[115]}), .b4_nUAi({
        b4_nUAi[784], b4_nUAi[783]}), .N_27(N_27_95), .N_25(N_25_95));
    b8_1LbcQDr1_x_252_0 b9_1LbcgKGIl (.mdiclink_reg({mdiclink_reg[124]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[252]}), .b4_nUAi({
        b4_nUAi[373], b4_nUAi[372]}), .N_27(N_27_43), .N_25(N_25_43));
    b8_1LbcQDr1_x_329_0 b8_1LbcgKEJ0 (.mdiclink_reg({mdiclink_reg[47]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[329]}), .b4_nUAi({
        b4_nUAi[142], b4_nUAi[141]}), .N_27(N_27_16), .N_25(N_25_16));
    b8_1LbcQDr1_x_257_0 b9_1LbcgKGSq (.mdiclink_reg({mdiclink_reg[119]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[257]}), .b4_nUAi({
        b4_nUAi[359], b4_nUAi[358], b4_nUAi[357]}), .b6_2ZTGIf({
        \b6_2ZTGIf[119] }));
    b8_1LbcQDr1_x_250_0 b9_1LbcgKGI5 (.mdiclink_reg({mdiclink_reg[126]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[250]}), .b4_nUAi({
        b4_nUAi[379], b4_nUAi[378]}), .N_27(N_27_45), .N_25(N_25_45));
    b8_1LbcQDr1_x_2_0 b9_1LbcgKeJl (.mdiclink_reg({mdiclink_reg[374]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[2]}), .b4_nUAi({
        b4_nUAi[1123], b4_nUAi[1122]}), .N_27(N_27_140), .N_25(
        N_25_140));
    b8_1LbcQDr1_x_245_0 b9_1LbcgKGqn (.mdiclink_reg({mdiclink_reg[131]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[245]}), .b4_nUAi({
        b4_nUAi[395], b4_nUAi[394], b4_nUAi[393]}), .b6_2ZTGIf({
        \b6_2ZTGIf[131] }));
    b8_1LbcQDr1_x_267_0 b9_1LbcgKGRq (.mdiclink_reg({mdiclink_reg[109]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[267]}), .b4_nUAi({
        b4_nUAi[328], b4_nUAi[327]}), .N_27(N_27_38), .N_25(N_25_38));
    b8_1LbcQDr1_x_106_0 b9_1LbcgKwJm (.mdiclink_reg({mdiclink_reg[270]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[106]}), .b4_nUAi({
        b4_nUAi[811], b4_nUAi[810]}), .N_27(N_27_99), .N_25(N_25_99));
    b8_1LbcQDr1_x_213_0 b9_1LbcgKGAV (.mdiclink_reg({mdiclink_reg[163]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[213]}), .b4_nUAi({
        b4_nUAi[491], b4_nUAi[490], b4_nUAi[489]}), .b6_2ZTGIf({
        \b6_2ZTGIf[163] }));
    b8_1LbcQDr1_x_135_0 b9_1LbcgKwQn0 (.mdiclink_reg({
        mdiclink_reg[241]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[135]}), 
        .b4_nUAi({b4_nUAi[725], b4_nUAi[724], b4_nUAi[723]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[241] }));
    b8_1LbcQDr1_x_258_0 b9_1LbcgKGSS (.mdiclink_reg({mdiclink_reg[118]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[258]}), .b4_nUAi({
        b4_nUAi[356], b4_nUAi[355], b4_nUAi[354]}), .b6_2ZTGIf({
        \b6_2ZTGIf[118] }));
    b8_1LbcQDr1_x_277_0 b8_1LbcgKJV (.mdiclink_reg({mdiclink_reg[99]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[277]}), .b4_nUAi({
        b4_nUAi[299], b4_nUAi[298], b4_nUAi[297]}), .b6_2ZTGIf({
        \b6_2ZTGIf[99] }));
    b8_1LbcQDr1_x_44_0 b9_1LbcgKeqd (.mdiclink_reg({mdiclink_reg[332]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[44]}), .b4_nUAi({
        b4_nUAi[997], b4_nUAi[996]}), .N_27(N_27_121), .N_25(N_25_121));
    b8_1LbcQDr1_x_341_0 b8_1LbcgKeU (.mdiclink_reg({mdiclink_reg[35]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[341]}), .b4_nUAi({
        b4_nUAi[107], b4_nUAi[106], b4_nUAi[105]}), .b6_2ZTGIf({
        \b6_2ZTGIf[35] }));
    b8_1LbcQDr1_x_147_0 b9_1LbcgKwIq (.mdiclink_reg({mdiclink_reg[229]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[147]}), .b4_nUAi({
        b4_nUAi[688], b4_nUAi[687]}), .N_27(N_27_83), .N_25(N_25_83));
    b8_1LbcQDr1_x_268_0 b9_1LbcgKGRS (.mdiclink_reg({mdiclink_reg[108]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[268]}), .b4_nUAi({
        b4_nUAi[325], b4_nUAi[324]}), .N_27(N_27_37), .N_25(N_25_37));
    b8_1LbcQDr1_x_6_0 b9_1LbcgKeJm (.mdiclink_reg({mdiclink_reg[370]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[6]}), .b4_nUAi({
        b4_nUAi[1111], b4_nUAi[1110]}), .N_27(N_27_138), .N_25(
        N_25_138));
    b8_1LbcQDr1_x_373_0 b7_1LbcgKe (.mdiclink_reg({mdiclink_reg[3]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[373]}), .b4_nUAi({
        b4_nUAi[11], b4_nUAi[10], b4_nUAi[9]}), .b6_2ZTGIf({
        \b6_2ZTGIf[3] }));
    b8_1LbcQDr1_x_259_0 b9_1LbcgKGSe (.mdiclink_reg({mdiclink_reg[117]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[259]}), .b4_nUAi({
        b4_nUAi[352], b4_nUAi[351]}), .N_27(N_27_41), .N_25(N_25_41));
    b8_1LbcQDr1_x_149_0 b9_1LbcgKwIe (.mdiclink_reg({mdiclink_reg[227]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[149]}), .b4_nUAi({
        b4_nUAi[683], b4_nUAi[682], b4_nUAi[681]}), .b6_2ZTGIf({
        \b6_2ZTGIf[227] }));
    b8_1LbcQDr1_x_233_0 b9_1LbcgKGQV0 (.mdiclink_reg({
        mdiclink_reg[143]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[233]}), 
        .b4_nUAi({b4_nUAi[430], b4_nUAi[429]}), .N_27(N_27_52), .N_25(
        N_25_52));
    b8_1LbcQDr1_x_269_0 b9_1LbcgKGRe (.mdiclink_reg({mdiclink_reg[107]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[269]}), .b4_nUAi({
        b4_nUAi[322], b4_nUAi[321]}), .N_27(N_27_36), .N_25(N_25_36));
    b8_1LbcQDr1_x_266_0 b9_1LbcgKGSm (.mdiclink_reg({mdiclink_reg[110]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[266]}), .b4_nUAi({
        b4_nUAi[331], b4_nUAi[330]}), .N_27(N_27_39), .N_25(N_25_39));
    b8_1LbcQDr1_x_276_0 b9_1LbcgKGRm (.mdiclink_reg({mdiclink_reg[100]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[276]}), .b4_nUAi({
        b4_nUAi[302], b4_nUAi[301], b4_nUAi[300]}), .b6_2ZTGIf({
        \b6_2ZTGIf[100] }));
    b8_1LbcQDr1_x_120_0 b9_1LbcgKwU5 (.mdiclink_reg({mdiclink_reg[256]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[120]}), .b4_nUAi({
        b4_nUAi[770], b4_nUAi[769], b4_nUAi[768]}), .b6_2ZTGIf({
        \b6_2ZTGIf[256] }));
    b8_1LbcQDr1_x_61_0 b9_1LbcgKeSp (.mdiclink_reg({mdiclink_reg[315]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[61]}), .b4_nUAi({
        b4_nUAi[946], b4_nUAi[945]}), .N_27(N_27_114), .N_25(N_25_114));
    b8_1LbcQDr1_x_295_0 b8_1LbcgKbS (.mdiclink_reg({mdiclink_reg[81]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[295]}), .b4_nUAi({
        b4_nUAi[245], b4_nUAi[244], b4_nUAi[243]}), .b6_2ZTGIf({
        \b6_2ZTGIf[81] }));
    b8_1LbcQDr1_x_71_0 b9_1LbcgKeRp (.mdiclink_reg({mdiclink_reg[305]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[71]}), .b4_nUAi({
        b4_nUAi[917], b4_nUAi[916], b4_nUAi[915]}), .b6_2ZTGIf({
        \b6_2ZTGIf[305] }));
    b8_1LbcQDr1_x_91_0 b9_1LbcgKwnp (.mdiclink_reg({mdiclink_reg[285]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[91]}), .b4_nUAi({
        b4_nUAi[856], b4_nUAi[855]}), .N_27(N_27_104), .N_25(N_25_104));
    b8_1LbcQDr1_x_296_0 b8_1LbcgKbR (.mdiclink_reg({mdiclink_reg[80]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[296]}), .b4_nUAi({
        b4_nUAi[242], b4_nUAi[241], b4_nUAi[240]}), .b6_2ZTGIf({
        \b6_2ZTGIf[80] }));
    b8_1LbcQDr1_x_194_0 b9_1LbcgKGnd (.mdiclink_reg({mdiclink_reg[182]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[194]}), .b4_nUAi({
        b4_nUAi[548], b4_nUAi[547], b4_nUAi[546]}), .b6_2ZTGIf({
        \b6_2ZTGIf[182] }));
    b8_1LbcQDr1_x_344_0 b8_1LbcgKeI (.mdiclink_reg({mdiclink_reg[32]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[344]}), .b4_nUAi({
        b4_nUAi[98], b4_nUAi[97], b4_nUAi[96]}), .b6_2ZTGIf({
        \b6_2ZTGIf[32] }));
    b8_1LbcQDr1_x_265_0 b9_1LbcgKGSn (.mdiclink_reg({mdiclink_reg[111]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[265]}), .b4_nUAi({
        b4_nUAi[334], b4_nUAi[333]}), .N_27(N_27_40), .N_25(N_25_40));
    b8_1LbcQDr1_x_37_0 b9_1LbcgKeqq (.mdiclink_reg({mdiclink_reg[339]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[37]}), .b4_nUAi({
        b4_nUAi[1019], b4_nUAi[1018], b4_nUAi[1017]}), .b6_2ZTGIf({
        \b6_2ZTGIf[339] }));
    b8_1LbcQDr1_x_353_0 b8_1LbcgKwq (.mdiclink_reg({mdiclink_reg[23]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[353]}), .b4_nUAi({
        b4_nUAi[71], b4_nUAi[70], b4_nUAi[69]}), .b6_2ZTGIf({
        \b6_2ZTGIf[23] }));
    b8_1LbcQDr1_x_313_0 b8_1LbcgKoq (.mdiclink_reg({mdiclink_reg[63]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[313]}), .b4_nUAi({
        b4_nUAi[190], b4_nUAi[189]}), .N_27(N_27_22), .N_25(N_25_22));
    b8_1LbcQDr1_x_275_0 b9_1LbcgKGRn (.mdiclink_reg({mdiclink_reg[101]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[275]}), .b4_nUAi({
        b4_nUAi[304], b4_nUAi[303]}), .N_27(N_27_35), .N_25(N_25_35));
    b8_1LbcQDr1_x_64_0 b9_1LbcgKeSd (.mdiclink_reg({mdiclink_reg[312]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[64]}), .b4_nUAi({
        b4_nUAi[938], b4_nUAi[937], b4_nUAi[936]}), .b6_2ZTGIf({
        \b6_2ZTGIf[312] }));
    b8_1LbcQDr1_x_81_0 b9_1LbcgKwVp (.mdiclink_reg({mdiclink_reg[295]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[81]}), .b4_nUAi({
        b4_nUAi[887], b4_nUAi[886], b4_nUAi[885]}), .b6_2ZTGIf({
        \b6_2ZTGIf[295] }));
    b8_1LbcQDr1_x_112_0 b9_1LbcgKwAl (.mdiclink_reg({mdiclink_reg[264]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[112]}), .b4_nUAi({
        b4_nUAi[794], b4_nUAi[793], b4_nUAi[792]}), .b6_2ZTGIf({
        \b6_2ZTGIf[264] }));
    b8_1LbcQDr1_x_74_0 b9_1LbcgKeRd (.mdiclink_reg({mdiclink_reg[302]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[74]}), .b4_nUAi({
        b4_nUAi[907], b4_nUAi[906]}), .N_27(N_27_111), .N_25(N_25_111));
    b8_1LbcQDr1_x_184_0 b9_1LbcgKGVd (.mdiclink_reg({mdiclink_reg[192]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[184]}), .b4_nUAi({
        b4_nUAi[578], b4_nUAi[577], b4_nUAi[576]}), .b6_2ZTGIf({
        \b6_2ZTGIf[192] }));
    b8_1LbcQDr1_x_145_0 b9_1LbcgKwqn (.mdiclink_reg({mdiclink_reg[231]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[145]}), .b4_nUAi({
        b4_nUAi[695], b4_nUAi[694], b4_nUAi[693]}), .b6_2ZTGIf({
        \b6_2ZTGIf[231] }));
    b8_1LbcQDr1_x_150_0 b9_1LbcgKwI5 (.mdiclink_reg({mdiclink_reg[226]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[150]}), .b4_nUAi({
        b4_nUAi[680], b4_nUAi[679], b4_nUAi[678]}), .b6_2ZTGIf({
        \b6_2ZTGIf[226] }));
    b8_1LbcQDr1_x_202_0 b9_1LbcgKGJl (.mdiclink_reg({mdiclink_reg[174]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[202]}), .b4_nUAi({
        b4_nUAi[523], b4_nUAi[522]}), .N_27(N_27_63), .N_25(N_25_63));
    b8_1LbcQDr1_x_132_0 b9_1LbcgKwQl0 (.mdiclink_reg({
        mdiclink_reg[244]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[132]}), 
        .b4_nUAi({b4_nUAi[734], b4_nUAi[733], b4_nUAi[732]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[244] }));
    b8_1LbcQDr1_x_191_0 b9_1LbcgKGnp (.mdiclink_reg({mdiclink_reg[185]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[191]}), .b4_nUAi({
        b4_nUAi[557], b4_nUAi[556], b4_nUAi[555]}), .b6_2ZTGIf({
        \b6_2ZTGIf[185] }));
    b8_1LbcQDr1_x_200_0 b9_1LbcgKGJ5 (.mdiclink_reg({mdiclink_reg[176]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[200]}), .b4_nUAi({
        b4_nUAi[530], b4_nUAi[529], b4_nUAi[528]}), .b6_2ZTGIf({
        \b6_2ZTGIf[176] }));
    b8_1LbcQDr1_x_10_0 b9_1LbcgKeA5 (.mdiclink_reg({mdiclink_reg[366]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[10]}), .b4_nUAi({
        b4_nUAi[1099], b4_nUAi[1098]}), .N_27(N_27_135), .N_25(
        N_25_135));
    b8_1LbcQDr1_x_243_0 b9_1LbcgKGqV (.mdiclink_reg({mdiclink_reg[133]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[243]}), .b4_nUAi({
        b4_nUAi[400], b4_nUAi[399]}), .N_27(N_27_47), .N_25(N_25_47));
    b8_1LbcQDr1_x_281_0 b8_1LbcgKJU (.mdiclink_reg({mdiclink_reg[95]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[281]}), .b4_nUAi({
        b4_nUAi[286], b4_nUAi[285]}), .N_27(N_27_34), .N_25(N_25_34));
    b8_1LbcQDr1_x_368_0 b7_1LbcgKb (.mdiclink_reg({mdiclink_reg[8]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[368]}), .b4_nUAi({
        b4_nUAi[26], b4_nUAi[25], b4_nUAi[24]}), .b6_2ZTGIf({
        \b6_2ZTGIf[8] }));
    b8_1LbcQDr1_x_97_0 b9_1LbcgKwJq (.mdiclink_reg({mdiclink_reg[279]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[97]}), .b4_nUAi({
        b4_nUAi[839], b4_nUAi[838], b4_nUAi[837]}), .b6_2ZTGIf({
        \b6_2ZTGIf[279] }));
    b8_1LbcQDr1_x_30_0 b9_1LbcgKeQ50 (.mdiclink_reg({mdiclink_reg[346]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[30]}), .b4_nUAi({
        b4_nUAi[1040], b4_nUAi[1039], b4_nUAi[1038]}), .b6_2ZTGIf({
        \b6_2ZTGIf[346] }));
    b8_1LbcQDr1_x_187_0 b9_1LbcgKGnq (.mdiclink_reg({mdiclink_reg[189]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[187]}), .b4_nUAi({
        b4_nUAi[568], b4_nUAi[567]}), .N_27(N_27_68), .N_25(N_25_68));
    b8_1LbcQDr1_x_181_0 b9_1LbcgKGVp (.mdiclink_reg({mdiclink_reg[195]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[181]}), .b4_nUAi({
        b4_nUAi[587], b4_nUAi[586], b4_nUAi[585]}), .b6_2ZTGIf({
        \b6_2ZTGIf[195] }));
    b8_1LbcQDr1_x_99_0 b9_1LbcgKwJe (.mdiclink_reg({mdiclink_reg[277]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[99]}), .b4_nUAi({
        b4_nUAi[832], b4_nUAi[831]}), .N_27(N_27_101), .N_25(N_25_101));
    b8_1LbcQDr1_x_57_0 b9_1LbcgKeSq (.mdiclink_reg({mdiclink_reg[319]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[57]}), .b4_nUAi({
        b4_nUAi[958], b4_nUAi[957]}), .N_27(N_27_118), .N_25(N_25_118));
    b8_1LbcQDr1_x_355_0 b8_1LbcgKwS (.mdiclink_reg({mdiclink_reg[21]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[355]}), .b4_nUAi({
        b4_nUAi[64], b4_nUAi[63]}), .N_27(N_27_5), .N_25(N_25_5));
    b8_1LbcQDr1_x_188_0 b9_1LbcgKGnS (.mdiclink_reg({mdiclink_reg[188]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[188]}), .b4_nUAi({
        b4_nUAi[565], b4_nUAi[564]}), .N_27(N_27_67), .N_25(N_25_67));
    b8_1LbcQDr1_x_315_0 b8_1LbcgKoS (.mdiclink_reg({mdiclink_reg[61]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[315]}), .b4_nUAi({
        b4_nUAi[184], b4_nUAi[183]}), .N_27(N_27_20), .N_25(N_25_20));
    b8_1LbcQDr1_x_67_0 b9_1LbcgKeRq (.mdiclink_reg({mdiclink_reg[309]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[67]}), .b4_nUAi({
        b4_nUAi[928], b4_nUAi[927]}), .N_27(N_27_113), .N_25(N_25_113));
    b8_1LbcQDr1_x_9_0 b9_1LbcgKeAe (.mdiclink_reg({mdiclink_reg[367]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[9]}), .b4_nUAi({
        b4_nUAi[1102], b4_nUAi[1101]}), .N_27(N_27_136), .N_25(
        N_25_136));
    b8_1LbcQDr1_x_356_0 b8_1LbcgKwR (.mdiclink_reg({mdiclink_reg[20]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[356]}), .b4_nUAi({
        b4_nUAi[62], b4_nUAi[61], b4_nUAi[60]}), .b6_2ZTGIf({
        \b6_2ZTGIf[20] }));
    b8_1LbcQDr1_x_23_0 b9_1LbcgKeUV (.mdiclink_reg({mdiclink_reg[353]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[23]}), .b4_nUAi({
        b4_nUAi[1061], b4_nUAi[1060], b4_nUAi[1059]}), .b6_2ZTGIf({
        \b6_2ZTGIf[353] }));
    b8_1LbcQDr1_x_316_0 b8_1LbcgKoR (.mdiclink_reg({mdiclink_reg[60]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[316]}), .b4_nUAi({
        b4_nUAi[181], b4_nUAi[180]}), .N_27(N_27_19), .N_25(N_25_19));
    b8_1LbcQDr1_x_189_0 b9_1LbcgKGne (.mdiclink_reg({mdiclink_reg[187]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[189]}), .b4_nUAi({
        b4_nUAi[562], b4_nUAi[561]}), .N_27(N_27_66), .N_25(N_25_66));
    b8_1LbcQDr1_x_177_0 b9_1LbcgKGVq (.mdiclink_reg({mdiclink_reg[199]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[177]}), .b4_nUAi({
        b4_nUAi[599], b4_nUAi[598], b4_nUAi[597]}), .b6_2ZTGIf({
        \b6_2ZTGIf[199] }));
    b8_1LbcQDr1_x_165_0 b9_1LbcgKwSn (.mdiclink_reg({mdiclink_reg[211]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[165]}), .b4_nUAi({
        b4_nUAi[635], b4_nUAi[634], b4_nUAi[633]}), .b6_2ZTGIf({
        \b6_2ZTGIf[211] }));
    b8_1LbcQDr1_x_29_0 b9_1LbcgKeQe0 (.mdiclink_reg({mdiclink_reg[347]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[29]}), .b4_nUAi({
        b4_nUAi[1042], b4_nUAi[1041]}), .N_27(N_27_126), .N_25(
        N_25_126));
    b8_1LbcQDr1_x_196_0 b9_1LbcgKGnm (.mdiclink_reg({mdiclink_reg[180]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[196]}), .b4_nUAi({
        b4_nUAi[542], b4_nUAi[541], b4_nUAi[540]}), .b6_2ZTGIf({
        \b6_2ZTGIf[180] }));
    b8_1LbcQDr1_x_114_0 b9_1LbcgKwAd (.mdiclink_reg({mdiclink_reg[262]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[114]}), .b4_nUAi({
        b4_nUAi[788], b4_nUAi[787], b4_nUAi[786]}), .b6_2ZTGIf({
        \b6_2ZTGIf[262] }));
    b8_1LbcQDr1_x_178_0 b9_1LbcgKGVS (.mdiclink_reg({mdiclink_reg[198]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[178]}), .b4_nUAi({
        b4_nUAi[596], b4_nUAi[595], b4_nUAi[594]}), .b6_2ZTGIf({
        \b6_2ZTGIf[198] }));
    b8_1LbcQDr1_x_284_0 b8_1LbcgKJI (.mdiclink_reg({mdiclink_reg[92]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[284]}), .b4_nUAi({
        b4_nUAi[277], b4_nUAi[276]}), .N_27(N_27_31), .N_25(N_25_31));
    b8_1LbcQDr1_x_175_0 b9_1LbcgKwRn (.mdiclink_reg({mdiclink_reg[201]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[175]}), .b4_nUAi({
        b4_nUAi[605], b4_nUAi[604], b4_nUAi[603]}), .b6_2ZTGIf({
        \b6_2ZTGIf[201] }));
    b8_1LbcQDr1_x_300_0 b8_1LbcgKxA (.mdiclink_reg({mdiclink_reg[76]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[300]}), .b4_nUAi({
        b4_nUAi[229], b4_nUAi[228]}), .N_27(N_27_25), .N_25(N_25_25));
    b8_1LbcQDr1_x_360_0 b8_1LbcgKGA (.mdiclink_reg({mdiclink_reg[16]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[360]}), .b4_nUAi({
        b4_nUAi[50], b4_nUAi[49], b4_nUAi[48]}), .b6_2ZTGIf({
        \b6_2ZTGIf[16] }));
    b8_1LbcQDr1_x_339_0 b8_1LbcgKeJ (.mdiclink_reg({mdiclink_reg[37]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[339]}), .b4_nUAi({
        b4_nUAi[112], b4_nUAi[111]}), .N_27(N_27_11), .N_25(N_25_11));
    b8_1LbcQDr1_x_179_0 b9_1LbcgKGVe (.mdiclink_reg({mdiclink_reg[197]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[179]}), .b4_nUAi({
        b4_nUAi[592], b4_nUAi[591]}), .N_27(N_27_71), .N_25(N_25_71));
    b8_1LbcQDr1_x_263_0 b9_1LbcgKGSV (.mdiclink_reg({mdiclink_reg[113]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[263]}), .b4_nUAi({
        b4_nUAi[341], b4_nUAi[340], b4_nUAi[339]}), .b6_2ZTGIf({
        \b6_2ZTGIf[113] }));
    b8_1LbcQDr1_x_288_0 b8_1LbcgKbn (.mdiclink_reg({mdiclink_reg[88]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[288]}), .b4_nUAi({
        b4_nUAi[266], b4_nUAi[265], b4_nUAi[264]}), .b6_2ZTGIf({
        \b6_2ZTGIf[88] }));
    b8_1LbcQDr1_x_134_0 b9_1LbcgKwQd0 (.mdiclink_reg({
        mdiclink_reg[242]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[134]}), 
        .b4_nUAi({b4_nUAi[728], b4_nUAi[727], b4_nUAi[726]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[242] }));
    b8_1LbcQDr1_x_273_0 b9_1LbcgKGRV (.mdiclink_reg({mdiclink_reg[103]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[273]}), .b4_nUAi({
        b4_nUAi[311], b4_nUAi[310], b4_nUAi[309]}), .b6_2ZTGIf({
        \b6_2ZTGIf[103] }));
    b8_1LbcQDr1_x_320_0 b8_1LbcgKIA (.mdiclink_reg({mdiclink_reg[56]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[320]}), .b4_nUAi({
        b4_nUAi[170], b4_nUAi[169], b4_nUAi[168]}), .b6_2ZTGIf({
        \b6_2ZTGIf[56] }));
    b8_1LbcQDr1_x_121_0 b9_1LbcgKwUp (.mdiclink_reg({mdiclink_reg[255]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[121]}), .b4_nUAi({
        b4_nUAi[766], b4_nUAi[765]}), .N_27(N_27_94), .N_25(N_25_94));
    b8_1LbcQDr1_x_142_0 b9_1LbcgKwql (.mdiclink_reg({mdiclink_reg[234]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[142]}), .b4_nUAi({
        b4_nUAi[704], b4_nUAi[703], b4_nUAi[702]}), .b6_2ZTGIf({
        \b6_2ZTGIf[234] }));
    b8_1LbcQDr1_x_186_0 b9_1LbcgKGVm (.mdiclink_reg({mdiclink_reg[190]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[186]}), .b4_nUAi({
        b4_nUAi[571], b4_nUAi[570]}), .N_27(N_27_69), .N_25(N_25_69));
    b8_1LbcQDr1_x_292_0 b8_1LbcgKbQ0 (.mdiclink_reg({mdiclink_reg[84]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[292]}), .b4_nUAi({
        b4_nUAi[254], b4_nUAi[253], b4_nUAi[252]}), .b6_2ZTGIf({
        \b6_2ZTGIf[84] }));
    b8_1LbcQDr1_x_224_0 b9_1LbcgKGUd (.mdiclink_reg({mdiclink_reg[152]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[224]}), .b4_nUAi({
        b4_nUAi[458], b4_nUAi[457], b4_nUAi[456]}), .b6_2ZTGIf({
        \b6_2ZTGIf[152] }));
    b8_1LbcQDr1_x_195_0 b9_1LbcgKGnn (.mdiclink_reg({mdiclink_reg[181]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[195]}), .b4_nUAi({
        b4_nUAi[544], b4_nUAi[543]}), .N_27(N_27_65), .N_25(N_25_65));
    b8_1LbcQDr1_x_53_0 b9_1LbcgKeIV (.mdiclink_reg({mdiclink_reg[323]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[53]}), .b4_nUAi({
        b4_nUAi[971], b4_nUAi[970], b4_nUAi[969]}), .b6_2ZTGIf({
        \b6_2ZTGIf[323] }));
    b8_1LbcQDr1_x_15_0 b9_1LbcgKeAn (.mdiclink_reg({mdiclink_reg[361]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[15]}), .b4_nUAi({
        b4_nUAi[1085], b4_nUAi[1084], b4_nUAi[1083]}), .b6_2ZTGIf({
        \b6_2ZTGIf[361] }));
    b8_1LbcQDr1_x_100_0 b9_1LbcgKwJ5 (.mdiclink_reg({mdiclink_reg[276]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[100]}), .b4_nUAi({
        b4_nUAi[830], b4_nUAi[829], b4_nUAi[828]}), .b6_2ZTGIf({
        \b6_2ZTGIf[276] }));
    b8_1LbcQDr1_x_40_0 b9_1LbcgKeq5 (.mdiclink_reg({mdiclink_reg[336]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[40]}), .b4_nUAi({
        b4_nUAi[1010], b4_nUAi[1009], b4_nUAi[1008]}), .b6_2ZTGIf({
        \b6_2ZTGIf[336] }));
    b8_1LbcQDr1_x_287_0 b8_1LbcgKbV (.mdiclink_reg({mdiclink_reg[89]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[287]}), .b4_nUAi({
        b4_nUAi[269], b4_nUAi[268], b4_nUAi[267]}), .b6_2ZTGIf({
        \b6_2ZTGIf[89] }));
    b8_1LbcQDr1_x_35_0 b9_1LbcgKeQn0 (.mdiclink_reg({mdiclink_reg[341]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[35]}), .b4_nUAi({
        b4_nUAi[1024], b4_nUAi[1023]}), .N_27(N_27_125), .N_25(
        N_25_125));
    b8_1LbcQDr1_x_185_0 b9_1LbcgKGVn (.mdiclink_reg({mdiclink_reg[191]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[185]}), .b4_nUAi({
        b4_nUAi[574], b4_nUAi[573]}), .N_27(N_27_70), .N_25(N_25_70));
    b8_1LbcQDr1_x_375_0 b7_1LbcgKG (.mdiclink_reg({mdiclink_reg[1]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[375]}), .b4_nUAi({b4_nUAi[5], 
        b4_nUAi[4], b4_nUAi[3]}), .b6_2ZTGIf({\b6_2ZTGIf[1] }));
    b8_1LbcQDr1_x_113_0 b9_1LbcgKwAV (.mdiclink_reg({mdiclink_reg[263]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[113]}), .b4_nUAi({
        b4_nUAi[791], b4_nUAi[790], b4_nUAi[789]}), .b6_2ZTGIf({
        \b6_2ZTGIf[263] }));
    b8_1LbcQDr1_x_221_0 b9_1LbcgKGUp (.mdiclink_reg({mdiclink_reg[155]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[221]}), .b4_nUAi({
        b4_nUAi[466], b4_nUAi[465]}), .N_27(N_27_54), .N_25(N_25_54));
    b8_1LbcQDr1_x_282_0 b8_1LbcgKJQ0 (.mdiclink_reg({mdiclink_reg[94]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[282]}), .b4_nUAi({
        b4_nUAi[283], b4_nUAi[282]}), .N_27(N_27_33), .N_25(N_25_33));
    b8_1LbcQDr1_x_151_0 b9_1LbcgKwIp (.mdiclink_reg({mdiclink_reg[225]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[151]}), .b4_nUAi({
        b4_nUAi[677], b4_nUAi[676], b4_nUAi[675]}), .b6_2ZTGIf({
        \b6_2ZTGIf[225] }));
    b8_1LbcQDr1_x_254_0 b9_1LbcgKGId (.mdiclink_reg({mdiclink_reg[122]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[254]}), .b4_nUAi({
        b4_nUAi[368], b4_nUAi[367], b4_nUAi[366]}), .b6_2ZTGIf({
        \b6_2ZTGIf[122] }));
    b8_1LbcQDr1_x_39_0 b9_1LbcgKeqe (.mdiclink_reg({mdiclink_reg[337]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[39]}), .b4_nUAi({
        b4_nUAi[1013], b4_nUAi[1012], b4_nUAi[1011]}), .b6_2ZTGIf({
        \b6_2ZTGIf[337] }));
    b8_1LbcQDr1_x_367_0 b7_1LbcgKJ (.mdiclink_reg({mdiclink_reg[9]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[367]}), .b4_nUAi({
        b4_nUAi[29], b4_nUAi[28], b4_nUAi[27]}), .b6_2ZTGIf({
        \b6_2ZTGIf[9] }));
    b8_1LbcQDr1_x_133_0 b9_1LbcgKwQV0 (.mdiclink_reg({
        mdiclink_reg[243]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[133]}), 
        .b4_nUAi({b4_nUAi[731], b4_nUAi[730], b4_nUAi[729]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[243] }));
    b8_1LbcQDr1_x_162_0 b9_1LbcgKwSl (.mdiclink_reg({mdiclink_reg[214]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[162]}), .b4_nUAi({
        b4_nUAi[644], b4_nUAi[643], b4_nUAi[642]}), .b6_2ZTGIf({
        \b6_2ZTGIf[214] }));
    b8_1LbcQDr1_x_217_0 b9_1LbcgKGUq (.mdiclink_reg({mdiclink_reg[159]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[217]}), .b4_nUAi({
        b4_nUAi[478], b4_nUAi[477]}), .N_27(N_27_58), .N_25(N_25_58));
    b8_1LbcQDr1_x_172_0 b9_1LbcgKwRl (.mdiclink_reg({mdiclink_reg[204]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[172]}), .b4_nUAi({
        b4_nUAi[613], b4_nUAi[612]}), .N_27(N_27_73), .N_25(N_25_73));
    b8_1LbcQDr1_x_348_0 b8_1LbcgKwn (.mdiclink_reg({mdiclink_reg[28]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[348]}), .b4_nUAi({
        b4_nUAi[85], b4_nUAi[84]}), .N_27(N_27_7), .N_25(N_25_7));
    b8_1LbcQDr1_x_144_0 b9_1LbcgKwqd (.mdiclink_reg({mdiclink_reg[232]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[144]}), .b4_nUAi({
        b4_nUAi[698], b4_nUAi[697], b4_nUAi[696]}), .b6_2ZTGIf({
        \b6_2ZTGIf[232] }));
    b8_1LbcQDr1_x_218_0 b9_1LbcgKGUS (.mdiclink_reg({mdiclink_reg[158]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[218]}), .b4_nUAi({
        b4_nUAi[475], b4_nUAi[474]}), .N_27(N_27_57), .N_25(N_25_57));
    b8_1LbcQDr1_x_308_0 b8_1LbcgKon (.mdiclink_reg({mdiclink_reg[68]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[308]}), .b4_nUAi({
        b4_nUAi[206], b4_nUAi[205], b4_nUAi[204]}), .b6_2ZTGIf({
        \b6_2ZTGIf[68] }));
    b8_1LbcQDr1_x_279_0 b8_1LbcgKJJ (.mdiclink_reg({mdiclink_reg[97]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[279]}), .b4_nUAi({
        b4_nUAi[293], b4_nUAi[292], b4_nUAi[291]}), .b6_2ZTGIf({
        \b6_2ZTGIf[97] }));
    b8_1LbcQDr1_x_60_0 b9_1LbcgKeS5 (.mdiclink_reg({mdiclink_reg[316]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[60]}), .b4_nUAi({
        b4_nUAi[949], b4_nUAi[948]}), .N_27(N_27_115), .N_25(N_25_115));
    b8_1LbcQDr1_x_303_0 b8_1LbcgKxq (.mdiclink_reg({mdiclink_reg[73]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[303]}), .b4_nUAi({
        b4_nUAi[221], b4_nUAi[220], b4_nUAi[219]}), .b6_2ZTGIf({
        \b6_2ZTGIf[73] }));
    b8_1LbcQDr1_x_363_0 b8_1LbcgKGq (.mdiclink_reg({mdiclink_reg[13]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[363]}), .b4_nUAi({
        b4_nUAi[40], b4_nUAi[39]}), .N_27(N_27_2), .N_25(N_25_2));
    b8_1LbcQDr1_x_108_0 b9_1LbcgKwAS (.mdiclink_reg({mdiclink_reg[268]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[108]}), .b4_nUAi({
        b4_nUAi[805], b4_nUAi[804]}), .N_27(N_27_97), .N_25(N_25_97));
    b8_1LbcQDr1_x_333_0 b8_1LbcgKEq0 (.mdiclink_reg({mdiclink_reg[43]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[333]}), .b4_nUAi({
        b4_nUAi[130], b4_nUAi[129]}), .N_27(N_27_12), .N_25(N_25_12));
    b8_1LbcQDr1_x_219_0 b9_1LbcgKGUe (.mdiclink_reg({mdiclink_reg[157]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[219]}), .b4_nUAi({
        b4_nUAi[472], b4_nUAi[471]}), .N_27(N_27_56), .N_25(N_25_56));
    b8_1LbcQDr1_x_70_0 b9_1LbcgKeR5 (.mdiclink_reg({mdiclink_reg[306]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[70]}), .b4_nUAi({
        b4_nUAi[920], b4_nUAi[919], b4_nUAi[918]}), .b6_2ZTGIf({
        \b6_2ZTGIf[306] }));
    b8_1LbcQDr1_x_251_0 b9_1LbcgKGIp (.mdiclink_reg({mdiclink_reg[125]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[251]}), .b4_nUAi({
        b4_nUAi[376], b4_nUAi[375]}), .N_27(N_27_44), .N_25(N_25_44));
    b8_1LbcQDr1_x_323_0 b8_1LbcgKIq (.mdiclink_reg({mdiclink_reg[53]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[323]}), .b4_nUAi({
        b4_nUAi[160], b4_nUAi[159]}), .N_27(N_27_17), .N_25(N_25_17));
    b8_1LbcQDr1_x_95_0 b9_1LbcgKwnn (.mdiclink_reg({mdiclink_reg[281]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[95]}), .b4_nUAi({
        b4_nUAi[845], b4_nUAi[844], b4_nUAi[843]}), .b6_2ZTGIf({
        \b6_2ZTGIf[281] }));
    b8_1LbcQDr1_x_347_0 b8_1LbcgKwV (.mdiclink_reg({mdiclink_reg[29]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[347]}), .b4_nUAi({
        b4_nUAi[88], b4_nUAi[87]}), .N_27(N_27_8), .N_25(N_25_8));
    b8_1LbcQDr1_x_226_0 b9_1LbcgKGUm (.mdiclink_reg({mdiclink_reg[150]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[226]}), .b4_nUAi({
        b4_nUAi[452], b4_nUAi[451], b4_nUAi[450]}), .b6_2ZTGIf({
        \b6_2ZTGIf[150] }));
    b8_1LbcQDr1_x_128_0 b9_1LbcgKwQS0 (.mdiclink_reg({
        mdiclink_reg[248]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[128]}), 
        .b4_nUAi({b4_nUAi[746], b4_nUAi[745], b4_nUAi[744]}), 
        .b6_2ZTGIf({\b6_2ZTGIf[248] }));
    b8_1LbcQDr1_x_307_0 b8_1LbcgKoV (.mdiclink_reg({mdiclink_reg[69]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[307]}), .b4_nUAi({
        b4_nUAi[208], b4_nUAi[207]}), .N_27(N_27_23), .N_25(N_25_23));
    b8_1LbcQDr1_x_330_0 b8_1LbcgKEA0 (.mdiclink_reg({mdiclink_reg[46]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[330]}), .b4_nUAi({
        b4_nUAi[139], b4_nUAi[138]}), .N_27(N_27_15), .N_25(N_25_15));
    b8_1LbcQDr1_x_12_0 b9_1LbcgKeAl (.mdiclink_reg({mdiclink_reg[364]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[12]}), .b4_nUAi({
        b4_nUAi[1093], b4_nUAi[1092]}), .N_27(N_27_133), .N_25(
        N_25_133));
    b8_1LbcQDr1_x_193_0 b9_1LbcgKGnV (.mdiclink_reg({mdiclink_reg[183]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[193]}), .b4_nUAi({
        b4_nUAi[551], b4_nUAi[550], b4_nUAi[549]}), .b6_2ZTGIf({
        \b6_2ZTGIf[183] }));
    b8_1LbcQDr1_x_45_0 b9_1LbcgKeqn (.mdiclink_reg({mdiclink_reg[331]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[45]}), .b4_nUAi({
        b4_nUAi[994], b4_nUAi[993]}), .N_27(N_27_120), .N_25(N_25_120));
    b8_1LbcQDr1_x_21_0 b9_1LbcgKeUp (.mdiclink_reg({mdiclink_reg[355]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[21]}), .b4_nUAi({
        b4_nUAi[1067], b4_nUAi[1066], b4_nUAi[1065]}), .b6_2ZTGIf({
        \b6_2ZTGIf[355] }));
    b8_1LbcQDr1_x_3_0 b9_1LbcgKeJV (.mdiclink_reg({mdiclink_reg[373]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[3]}), .b4_nUAi({
        b4_nUAi[1121], b4_nUAi[1120], b4_nUAi[1119]}), .b6_2ZTGIf({
        \b6_2ZTGIf[373] }));
    b8_1LbcQDr1_x_116_0 b9_1LbcgKwAm (.mdiclink_reg({mdiclink_reg[260]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[116]}), .b4_nUAi({
        b4_nUAi[782], b4_nUAi[781], b4_nUAi[780]}), .b6_2ZTGIf({
        \b6_2ZTGIf[260] }));
    b8_1LbcQDr1_x_247_0 b9_1LbcgKGIq (.mdiclink_reg({mdiclink_reg[129]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[247]}), .b4_nUAi({
        b4_nUAi[389], b4_nUAi[388], b4_nUAi[387]}), .b6_2ZTGIf({
        \b6_2ZTGIf[129] }));
    b8_1LbcQDr1_x_59_0 b9_1LbcgKeSe (.mdiclink_reg({mdiclink_reg[317]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[59]}), .b4_nUAi({
        b4_nUAi[952], b4_nUAi[951]}), .N_27(N_27_116), .N_25(N_25_116));
    b8_1LbcQDr1_x_291_0 b8_1LbcgKbU (.mdiclink_reg({mdiclink_reg[85]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[291]}), .b4_nUAi({
        b4_nUAi[256], b4_nUAi[255]}), .N_27(N_27_29), .N_25(N_25_29));
    
endmodule


module b7_PfFzrNY_x_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       IICE_comm2iice,
       b11_PSyil9s_FMZ,
       BW_clk_c,
       b7_PSyi3wy,
       b4_PLyF,
       b8_PSyiBgYG
    );
input  [376:0] mdiclink_reg;
input  [376:0] b11_OFWNT9L_8tZ;
input  [11:10] IICE_comm2iice;
output b11_PSyil9s_FMZ;
input  BW_clk_c;
output b7_PSyi3wy;
input  b4_PLyF;
input  b8_PSyiBgYG;

    wire VCC_net_1, \b11_uUT0JC4gFrY[1] , GND_net_1, \b4_nUAi[0] , 
        \b4_nUAi[1] , \b4_nUAi[2] , \b4_nUAi[3] , \b4_nUAi[4] , 
        \b4_nUAi[5] , \b4_nUAi[6] , \b4_nUAi[7] , \b4_nUAi[8] , 
        \b4_nUAi[9] , \b4_nUAi[10] , \b4_nUAi[11] , \b4_nUAi[12] , 
        \b4_nUAi[13] , \b4_nUAi[14] , \b4_nUAi[15] , \b4_nUAi[16] , 
        \b4_nUAi[17] , \b4_nUAi[18] , \b4_nUAi[19] , \b4_nUAi[20] , 
        \b4_nUAi[21] , \b4_nUAi[22] , \b4_nUAi[23] , \b4_nUAi[24] , 
        \b4_nUAi[25] , \b4_nUAi[26] , \b4_nUAi[27] , \b4_nUAi[28] , 
        \b4_nUAi[29] , \b4_nUAi[30] , \b4_nUAi[31] , \b4_nUAi[32] , 
        \b4_nUAi[33] , \b4_nUAi[34] , \b4_nUAi[35] , \b4_nUAi[36] , 
        \b4_nUAi[37] , \b4_nUAi[38] , \b4_nUAi[39] , \b4_nUAi[40] , 
        \b4_nUAi[41] , \b4_nUAi[42] , \b4_nUAi[43] , \b4_nUAi[44] , 
        \b4_nUAi[45] , \b4_nUAi[46] , \b4_nUAi[47] , \b4_nUAi[48] , 
        \b4_nUAi[49] , \b4_nUAi[50] , \b4_nUAi[51] , \b4_nUAi[52] , 
        \b4_nUAi[53] , \b4_nUAi[54] , \b4_nUAi[55] , \b4_nUAi[56] , 
        \b4_nUAi[57] , \b4_nUAi[58] , \b4_nUAi[59] , \b4_nUAi[60] , 
        \b4_nUAi[61] , \b4_nUAi[62] , \b4_nUAi[63] , \b4_nUAi[64] , 
        \b4_nUAi[65] , \b4_nUAi[66] , \b4_nUAi[67] , \b4_nUAi[68] , 
        \b4_nUAi[69] , \b4_nUAi[70] , \b4_nUAi[71] , \b4_nUAi[72] , 
        \b4_nUAi[73] , \b4_nUAi[74] , \b4_nUAi[75] , \b4_nUAi[76] , 
        \b4_nUAi[77] , \b4_nUAi[78] , \b4_nUAi[79] , \b4_nUAi[80] , 
        \b4_nUAi[81] , \b4_nUAi[82] , \b4_nUAi[83] , \b4_nUAi[84] , 
        \b4_nUAi[85] , \b4_nUAi[86] , \b4_nUAi[87] , \b4_nUAi[88] , 
        \b4_nUAi[89] , \b4_nUAi[90] , \b4_nUAi[91] , \b4_nUAi[92] , 
        \b4_nUAi[93] , \b4_nUAi[94] , \b4_nUAi[95] , \b4_nUAi[96] , 
        \b4_nUAi[97] , \b4_nUAi[98] , \b4_nUAi[99] , \b4_nUAi[100] , 
        \b4_nUAi[101] , \b4_nUAi[102] , \b4_nUAi[103] , \b4_nUAi[104] , 
        \b4_nUAi[105] , \b4_nUAi[106] , \b4_nUAi[107] , \b4_nUAi[108] , 
        \b4_nUAi[109] , \b4_nUAi[110] , \b4_nUAi[111] , \b4_nUAi[112] , 
        \b4_nUAi[113] , \b4_nUAi[114] , \b4_nUAi[115] , \b4_nUAi[116] , 
        \b4_nUAi[117] , \b4_nUAi[118] , \b4_nUAi[119] , \b4_nUAi[120] , 
        \b4_nUAi[121] , \b4_nUAi[122] , \b4_nUAi[123] , \b4_nUAi[124] , 
        \b4_nUAi[125] , \b4_nUAi[126] , \b4_nUAi[127] , \b4_nUAi[128] , 
        \b4_nUAi[129] , \b4_nUAi[130] , \b4_nUAi[131] , \b4_nUAi[132] , 
        \b4_nUAi[133] , \b4_nUAi[134] , \b4_nUAi[135] , \b4_nUAi[136] , 
        \b4_nUAi[137] , \b4_nUAi[138] , \b4_nUAi[139] , \b4_nUAi[140] , 
        \b4_nUAi[141] , \b4_nUAi[142] , \b4_nUAi[143] , \b4_nUAi[144] , 
        \b4_nUAi[145] , \b4_nUAi[146] , \b4_nUAi[147] , \b4_nUAi[148] , 
        \b4_nUAi[149] , \b4_nUAi[150] , \b4_nUAi[151] , \b4_nUAi[152] , 
        \b4_nUAi[153] , \b4_nUAi[154] , \b4_nUAi[155] , \b4_nUAi[156] , 
        \b4_nUAi[157] , \b4_nUAi[158] , \b4_nUAi[159] , \b4_nUAi[160] , 
        \b4_nUAi[161] , \b4_nUAi[162] , \b4_nUAi[163] , \b4_nUAi[164] , 
        \b4_nUAi[165] , \b4_nUAi[166] , \b4_nUAi[167] , \b4_nUAi[168] , 
        \b4_nUAi[169] , \b4_nUAi[170] , \b4_nUAi[171] , \b4_nUAi[172] , 
        \b4_nUAi[173] , \b4_nUAi[174] , \b4_nUAi[175] , \b4_nUAi[176] , 
        \b4_nUAi[177] , \b4_nUAi[178] , \b4_nUAi[179] , \b4_nUAi[180] , 
        \b4_nUAi[181] , \b4_nUAi[182] , \b4_nUAi[183] , \b4_nUAi[184] , 
        \b4_nUAi[185] , \b4_nUAi[186] , \b4_nUAi[187] , \b4_nUAi[188] , 
        \b4_nUAi[189] , \b4_nUAi[190] , \b4_nUAi[191] , \b4_nUAi[192] , 
        \b4_nUAi[193] , \b4_nUAi[194] , \b4_nUAi[195] , \b4_nUAi[196] , 
        \b4_nUAi[197] , \b4_nUAi[198] , \b4_nUAi[199] , \b4_nUAi[200] , 
        \b4_nUAi[201] , \b4_nUAi[202] , \b4_nUAi[203] , \b4_nUAi[204] , 
        \b4_nUAi[205] , \b4_nUAi[206] , \b4_nUAi[207] , \b4_nUAi[208] , 
        \b4_nUAi[209] , \b4_nUAi[210] , \b4_nUAi[211] , \b4_nUAi[212] , 
        \b4_nUAi[213] , \b4_nUAi[214] , \b4_nUAi[215] , \b4_nUAi[216] , 
        \b4_nUAi[217] , \b4_nUAi[218] , \b4_nUAi[219] , \b4_nUAi[220] , 
        \b4_nUAi[221] , \b4_nUAi[222] , \b4_nUAi[223] , \b4_nUAi[224] , 
        \b4_nUAi[225] , \b4_nUAi[226] , \b4_nUAi[227] , \b4_nUAi[228] , 
        \b4_nUAi[229] , \b4_nUAi[230] , \b4_nUAi[231] , \b4_nUAi[232] , 
        \b4_nUAi[233] , \b4_nUAi[234] , \b4_nUAi[235] , \b4_nUAi[236] , 
        \b4_nUAi[237] , \b4_nUAi[238] , \b4_nUAi[239] , \b4_nUAi[240] , 
        \b4_nUAi[241] , \b4_nUAi[242] , \b4_nUAi[243] , \b4_nUAi[244] , 
        \b4_nUAi[245] , \b4_nUAi[246] , \b4_nUAi[247] , \b4_nUAi[248] , 
        \b4_nUAi[249] , \b4_nUAi[250] , \b4_nUAi[251] , \b4_nUAi[252] , 
        \b4_nUAi[253] , \b4_nUAi[254] , \b4_nUAi[255] , \b4_nUAi[256] , 
        \b4_nUAi[257] , \b4_nUAi[258] , \b4_nUAi[259] , \b4_nUAi[260] , 
        \b4_nUAi[261] , \b4_nUAi[262] , \b4_nUAi[263] , \b4_nUAi[264] , 
        \b4_nUAi[265] , \b4_nUAi[266] , \b4_nUAi[267] , \b4_nUAi[268] , 
        \b4_nUAi[269] , \b4_nUAi[270] , \b4_nUAi[271] , \b4_nUAi[272] , 
        \b4_nUAi[273] , \b4_nUAi[274] , \b4_nUAi[275] , \b4_nUAi[276] , 
        \b4_nUAi[277] , \b4_nUAi[278] , \b4_nUAi[279] , \b4_nUAi[280] , 
        \b4_nUAi[281] , \b4_nUAi[282] , \b4_nUAi[283] , \b4_nUAi[284] , 
        \b4_nUAi[285] , \b4_nUAi[286] , \b4_nUAi[287] , \b4_nUAi[288] , 
        \b4_nUAi[289] , \b4_nUAi[290] , \b4_nUAi[291] , \b4_nUAi[292] , 
        \b4_nUAi[293] , \b4_nUAi[294] , \b4_nUAi[295] , \b4_nUAi[296] , 
        \b4_nUAi[297] , \b4_nUAi[298] , \b4_nUAi[299] , \b4_nUAi[300] , 
        \b4_nUAi[301] , \b4_nUAi[302] , \b4_nUAi[303] , \b4_nUAi[304] , 
        \b4_nUAi[305] , \b4_nUAi[306] , \b4_nUAi[307] , \b4_nUAi[308] , 
        \b4_nUAi[309] , \b4_nUAi[310] , \b4_nUAi[311] , \b4_nUAi[312] , 
        \b4_nUAi[313] , \b4_nUAi[314] , \b4_nUAi[315] , \b4_nUAi[316] , 
        \b4_nUAi[317] , \b4_nUAi[318] , \b4_nUAi[319] , \b4_nUAi[320] , 
        \b4_nUAi[321] , \b4_nUAi[322] , \b4_nUAi[323] , \b4_nUAi[324] , 
        \b4_nUAi[325] , \b4_nUAi[326] , \b4_nUAi[327] , \b4_nUAi[328] , 
        \b4_nUAi[329] , \b4_nUAi[330] , \b4_nUAi[331] , \b4_nUAi[332] , 
        \b4_nUAi[333] , \b4_nUAi[334] , \b4_nUAi[335] , \b4_nUAi[336] , 
        \b4_nUAi[337] , \b4_nUAi[338] , \b4_nUAi[339] , \b4_nUAi[340] , 
        \b4_nUAi[341] , \b4_nUAi[342] , \b4_nUAi[343] , \b4_nUAi[344] , 
        \b4_nUAi[345] , \b4_nUAi[346] , \b4_nUAi[347] , \b4_nUAi[348] , 
        \b4_nUAi[349] , \b4_nUAi[350] , \b4_nUAi[351] , \b4_nUAi[352] , 
        \b4_nUAi[353] , \b4_nUAi[354] , \b4_nUAi[355] , \b4_nUAi[356] , 
        \b4_nUAi[357] , \b4_nUAi[358] , \b4_nUAi[359] , \b4_nUAi[360] , 
        \b4_nUAi[361] , \b4_nUAi[362] , \b4_nUAi[363] , \b4_nUAi[364] , 
        \b4_nUAi[365] , \b4_nUAi[366] , \b4_nUAi[367] , \b4_nUAi[368] , 
        \b4_nUAi[369] , \b4_nUAi[370] , \b4_nUAi[371] , \b4_nUAi[372] , 
        \b4_nUAi[373] , \b4_nUAi[374] , \b4_nUAi[375] , \b4_nUAi[376] , 
        \b4_nUAi[377] , \b4_nUAi[378] , \b4_nUAi[379] , \b4_nUAi[380] , 
        \b4_nUAi[381] , \b4_nUAi[382] , \b4_nUAi[383] , \b4_nUAi[384] , 
        \b4_nUAi[385] , \b4_nUAi[386] , \b4_nUAi[387] , \b4_nUAi[388] , 
        \b4_nUAi[389] , \b4_nUAi[390] , \b4_nUAi[391] , \b4_nUAi[392] , 
        \b4_nUAi[393] , \b4_nUAi[394] , \b4_nUAi[395] , \b4_nUAi[396] , 
        \b4_nUAi[397] , \b4_nUAi[398] , \b4_nUAi[399] , \b4_nUAi[400] , 
        \b4_nUAi[401] , \b4_nUAi[402] , \b4_nUAi[403] , \b4_nUAi[404] , 
        \b4_nUAi[405] , \b4_nUAi[406] , \b4_nUAi[407] , \b4_nUAi[408] , 
        \b4_nUAi[409] , \b4_nUAi[410] , \b4_nUAi[411] , \b4_nUAi[412] , 
        \b4_nUAi[413] , \b4_nUAi[414] , \b4_nUAi[415] , \b4_nUAi[416] , 
        \b4_nUAi[417] , \b4_nUAi[418] , \b4_nUAi[419] , \b4_nUAi[420] , 
        \b4_nUAi[421] , \b4_nUAi[422] , \b4_nUAi[423] , \b4_nUAi[424] , 
        \b4_nUAi[425] , \b4_nUAi[426] , \b4_nUAi[427] , \b4_nUAi[428] , 
        \b4_nUAi[429] , \b4_nUAi[430] , \b4_nUAi[431] , \b4_nUAi[432] , 
        \b4_nUAi[433] , \b4_nUAi[434] , \b4_nUAi[435] , \b4_nUAi[436] , 
        \b4_nUAi[437] , \b4_nUAi[438] , \b4_nUAi[439] , \b4_nUAi[440] , 
        \b4_nUAi[441] , \b4_nUAi[442] , \b4_nUAi[443] , \b4_nUAi[444] , 
        \b4_nUAi[445] , \b4_nUAi[446] , \b4_nUAi[447] , \b4_nUAi[448] , 
        \b4_nUAi[449] , \b4_nUAi[450] , \b4_nUAi[451] , \b4_nUAi[452] , 
        \b4_nUAi[453] , \b4_nUAi[454] , \b4_nUAi[455] , \b4_nUAi[456] , 
        \b4_nUAi[457] , \b4_nUAi[458] , \b4_nUAi[459] , \b4_nUAi[460] , 
        \b4_nUAi[461] , \b4_nUAi[462] , \b4_nUAi[463] , \b4_nUAi[464] , 
        \b4_nUAi[465] , \b4_nUAi[466] , \b4_nUAi[467] , \b4_nUAi[468] , 
        \b4_nUAi[469] , \b4_nUAi[470] , \b4_nUAi[471] , \b4_nUAi[472] , 
        \b4_nUAi[473] , \b4_nUAi[474] , \b4_nUAi[475] , \b4_nUAi[476] , 
        \b4_nUAi[477] , \b4_nUAi[478] , \b4_nUAi[479] , \b4_nUAi[480] , 
        \b4_nUAi[481] , \b4_nUAi[482] , \b4_nUAi[483] , \b4_nUAi[484] , 
        \b4_nUAi[485] , \b4_nUAi[486] , \b4_nUAi[487] , \b4_nUAi[488] , 
        \b4_nUAi[489] , \b4_nUAi[490] , \b4_nUAi[491] , \b4_nUAi[492] , 
        \b4_nUAi[493] , \b4_nUAi[494] , \b4_nUAi[495] , \b4_nUAi[496] , 
        \b4_nUAi[497] , \b4_nUAi[498] , \b4_nUAi[499] , \b4_nUAi[500] , 
        \b4_nUAi[501] , \b4_nUAi[502] , \b4_nUAi[503] , \b4_nUAi[504] , 
        \b4_nUAi[505] , \b4_nUAi[506] , \b4_nUAi[507] , \b4_nUAi[508] , 
        \b4_nUAi[509] , \b4_nUAi[510] , \b4_nUAi[511] , \b4_nUAi[512] , 
        \b4_nUAi[513] , \b4_nUAi[514] , \b4_nUAi[515] , \b4_nUAi[516] , 
        \b4_nUAi[517] , \b4_nUAi[518] , \b4_nUAi[519] , \b4_nUAi[520] , 
        \b4_nUAi[521] , \b4_nUAi[522] , \b4_nUAi[523] , \b4_nUAi[524] , 
        \b4_nUAi[525] , \b4_nUAi[526] , \b4_nUAi[527] , \b4_nUAi[528] , 
        \b4_nUAi[529] , \b4_nUAi[530] , \b4_nUAi[531] , \b4_nUAi[532] , 
        \b4_nUAi[533] , \b4_nUAi[534] , \b4_nUAi[535] , \b4_nUAi[536] , 
        \b4_nUAi[537] , \b4_nUAi[538] , \b4_nUAi[539] , \b4_nUAi[540] , 
        \b4_nUAi[541] , \b4_nUAi[542] , \b4_nUAi[543] , \b4_nUAi[544] , 
        \b4_nUAi[545] , \b4_nUAi[546] , \b4_nUAi[547] , \b4_nUAi[548] , 
        \b4_nUAi[549] , \b4_nUAi[550] , \b4_nUAi[551] , \b4_nUAi[552] , 
        \b4_nUAi[553] , \b4_nUAi[554] , \b4_nUAi[555] , \b4_nUAi[556] , 
        \b4_nUAi[557] , \b4_nUAi[558] , \b4_nUAi[559] , \b4_nUAi[560] , 
        \b4_nUAi[561] , \b4_nUAi[562] , \b4_nUAi[563] , \b4_nUAi[564] , 
        \b4_nUAi[565] , \b4_nUAi[566] , \b4_nUAi[567] , \b4_nUAi[568] , 
        \b4_nUAi[569] , \b4_nUAi[570] , \b4_nUAi[571] , \b4_nUAi[572] , 
        \b4_nUAi[573] , \b4_nUAi[574] , \b4_nUAi[575] , \b4_nUAi[576] , 
        \b4_nUAi[577] , \b4_nUAi[578] , \b4_nUAi[579] , \b4_nUAi[580] , 
        \b4_nUAi[581] , \b4_nUAi[582] , \b4_nUAi[583] , \b4_nUAi[584] , 
        \b4_nUAi[585] , \b4_nUAi[586] , \b4_nUAi[587] , \b4_nUAi[588] , 
        \b4_nUAi[589] , \b4_nUAi[590] , \b4_nUAi[591] , \b4_nUAi[592] , 
        \b4_nUAi[593] , \b4_nUAi[594] , \b4_nUAi[595] , \b4_nUAi[596] , 
        \b4_nUAi[597] , \b4_nUAi[598] , \b4_nUAi[599] , \b4_nUAi[600] , 
        \b4_nUAi[601] , \b4_nUAi[602] , \b4_nUAi[603] , \b4_nUAi[604] , 
        \b4_nUAi[605] , \b4_nUAi[606] , \b4_nUAi[607] , \b4_nUAi[608] , 
        \b4_nUAi[609] , \b4_nUAi[610] , \b4_nUAi[611] , \b4_nUAi[612] , 
        \b4_nUAi[613] , \b4_nUAi[614] , \b4_nUAi[615] , \b4_nUAi[616] , 
        \b4_nUAi[617] , \b4_nUAi[618] , \b4_nUAi[619] , \b4_nUAi[620] , 
        \b4_nUAi[621] , \b4_nUAi[622] , \b4_nUAi[623] , \b4_nUAi[624] , 
        \b4_nUAi[625] , \b4_nUAi[626] , \b4_nUAi[627] , \b4_nUAi[628] , 
        \b4_nUAi[629] , \b4_nUAi[630] , \b4_nUAi[631] , \b4_nUAi[632] , 
        \b4_nUAi[633] , \b4_nUAi[634] , \b4_nUAi[635] , \b4_nUAi[636] , 
        \b4_nUAi[637] , \b4_nUAi[638] , \b4_nUAi[639] , \b4_nUAi[640] , 
        \b4_nUAi[641] , \b4_nUAi[642] , \b4_nUAi[643] , \b4_nUAi[644] , 
        \b4_nUAi[645] , \b4_nUAi[646] , \b4_nUAi[647] , \b4_nUAi[648] , 
        \b4_nUAi[649] , \b4_nUAi[650] , \b4_nUAi[651] , \b4_nUAi[652] , 
        \b4_nUAi[653] , \b4_nUAi[654] , \b4_nUAi[655] , \b4_nUAi[656] , 
        \b4_nUAi[657] , \b4_nUAi[658] , \b4_nUAi[659] , \b4_nUAi[660] , 
        \b4_nUAi[661] , \b4_nUAi[662] , \b4_nUAi[663] , \b4_nUAi[664] , 
        \b4_nUAi[665] , \b4_nUAi[666] , \b4_nUAi[667] , \b4_nUAi[668] , 
        \b4_nUAi[669] , \b4_nUAi[670] , \b4_nUAi[671] , \b4_nUAi[672] , 
        \b4_nUAi[673] , \b4_nUAi[674] , \b4_nUAi[675] , \b4_nUAi[676] , 
        \b4_nUAi[677] , \b4_nUAi[678] , \b4_nUAi[679] , \b4_nUAi[680] , 
        \b4_nUAi[681] , \b4_nUAi[682] , \b4_nUAi[683] , \b4_nUAi[684] , 
        \b4_nUAi[685] , \b4_nUAi[686] , \b4_nUAi[687] , \b4_nUAi[688] , 
        \b4_nUAi[689] , \b4_nUAi[690] , \b4_nUAi[691] , \b4_nUAi[692] , 
        \b4_nUAi[693] , \b4_nUAi[694] , \b4_nUAi[695] , \b4_nUAi[696] , 
        \b4_nUAi[697] , \b4_nUAi[698] , \b4_nUAi[699] , \b4_nUAi[700] , 
        \b4_nUAi[701] , \b4_nUAi[702] , \b4_nUAi[703] , \b4_nUAi[704] , 
        \b4_nUAi[705] , \b4_nUAi[706] , \b4_nUAi[707] , \b4_nUAi[708] , 
        \b4_nUAi[709] , \b4_nUAi[710] , \b4_nUAi[711] , \b4_nUAi[712] , 
        \b4_nUAi[713] , \b4_nUAi[714] , \b4_nUAi[715] , \b4_nUAi[716] , 
        \b4_nUAi[717] , \b4_nUAi[718] , \b4_nUAi[719] , \b4_nUAi[720] , 
        \b4_nUAi[721] , \b4_nUAi[722] , \b4_nUAi[723] , \b4_nUAi[724] , 
        \b4_nUAi[725] , \b4_nUAi[726] , \b4_nUAi[727] , \b4_nUAi[728] , 
        \b4_nUAi[729] , \b4_nUAi[730] , \b4_nUAi[731] , \b4_nUAi[732] , 
        \b4_nUAi[733] , \b4_nUAi[734] , \b4_nUAi[735] , \b4_nUAi[736] , 
        \b4_nUAi[737] , \b4_nUAi[738] , \b4_nUAi[739] , \b4_nUAi[740] , 
        \b4_nUAi[741] , \b4_nUAi[742] , \b4_nUAi[743] , \b4_nUAi[744] , 
        \b4_nUAi[745] , \b4_nUAi[746] , \b4_nUAi[747] , \b4_nUAi[748] , 
        \b4_nUAi[749] , \b4_nUAi[750] , \b4_nUAi[751] , \b4_nUAi[752] , 
        \b4_nUAi[753] , \b4_nUAi[754] , \b4_nUAi[755] , \b4_nUAi[756] , 
        \b4_nUAi[757] , \b4_nUAi[758] , \b4_nUAi[759] , \b4_nUAi[760] , 
        \b4_nUAi[761] , \b4_nUAi[762] , \b4_nUAi[763] , \b4_nUAi[764] , 
        \b4_nUAi[765] , \b4_nUAi[766] , \b4_nUAi[767] , \b4_nUAi[768] , 
        \b4_nUAi[769] , \b4_nUAi[770] , \b4_nUAi[771] , \b4_nUAi[772] , 
        \b4_nUAi[773] , \b4_nUAi[774] , \b4_nUAi[775] , \b4_nUAi[776] , 
        \b4_nUAi[777] , \b4_nUAi[778] , \b4_nUAi[779] , \b4_nUAi[780] , 
        \b4_nUAi[781] , \b4_nUAi[782] , \b4_nUAi[783] , \b4_nUAi[784] , 
        \b4_nUAi[785] , \b4_nUAi[786] , \b4_nUAi[787] , \b4_nUAi[788] , 
        \b4_nUAi[789] , \b4_nUAi[790] , \b4_nUAi[791] , \b4_nUAi[792] , 
        \b4_nUAi[793] , \b4_nUAi[794] , \b4_nUAi[795] , \b4_nUAi[796] , 
        \b4_nUAi[797] , \b4_nUAi[798] , \b4_nUAi[799] , \b4_nUAi[800] , 
        \b4_nUAi[801] , \b4_nUAi[802] , \b4_nUAi[803] , \b4_nUAi[804] , 
        \b4_nUAi[805] , \b4_nUAi[806] , \b4_nUAi[807] , \b4_nUAi[808] , 
        \b4_nUAi[809] , \b4_nUAi[810] , \b4_nUAi[811] , \b4_nUAi[812] , 
        \b4_nUAi[813] , \b4_nUAi[814] , \b4_nUAi[815] , \b4_nUAi[816] , 
        \b4_nUAi[817] , \b4_nUAi[818] , \b4_nUAi[819] , \b4_nUAi[820] , 
        \b4_nUAi[821] , \b4_nUAi[822] , \b4_nUAi[823] , \b4_nUAi[824] , 
        \b4_nUAi[825] , \b4_nUAi[826] , \b4_nUAi[827] , \b4_nUAi[828] , 
        \b4_nUAi[829] , \b4_nUAi[830] , \b4_nUAi[831] , \b4_nUAi[832] , 
        \b4_nUAi[833] , \b4_nUAi[834] , \b4_nUAi[835] , \b4_nUAi[836] , 
        \b4_nUAi[837] , \b4_nUAi[838] , \b4_nUAi[839] , \b4_nUAi[840] , 
        \b4_nUAi[841] , \b4_nUAi[842] , \b4_nUAi[843] , \b4_nUAi[844] , 
        \b4_nUAi[845] , \b4_nUAi[846] , \b4_nUAi[847] , \b4_nUAi[848] , 
        \b4_nUAi[849] , \b4_nUAi[850] , \b4_nUAi[851] , \b4_nUAi[852] , 
        \b4_nUAi[853] , \b4_nUAi[854] , \b4_nUAi[855] , \b4_nUAi[856] , 
        \b4_nUAi[857] , \b4_nUAi[858] , \b4_nUAi[859] , \b4_nUAi[860] , 
        \b4_nUAi[861] , \b4_nUAi[862] , \b4_nUAi[863] , \b4_nUAi[864] , 
        \b4_nUAi[865] , \b4_nUAi[866] , \b4_nUAi[867] , \b4_nUAi[868] , 
        \b4_nUAi[869] , \b4_nUAi[870] , \b4_nUAi[871] , \b4_nUAi[872] , 
        \b4_nUAi[873] , \b4_nUAi[874] , \b4_nUAi[875] , \b4_nUAi[876] , 
        \b4_nUAi[877] , \b4_nUAi[878] , \b4_nUAi[879] , \b4_nUAi[880] , 
        \b4_nUAi[881] , \b4_nUAi[882] , \b4_nUAi[883] , \b4_nUAi[884] , 
        \b4_nUAi[885] , \b4_nUAi[886] , \b4_nUAi[887] , \b4_nUAi[888] , 
        \b4_nUAi[889] , \b4_nUAi[890] , \b4_nUAi[891] , \b4_nUAi[892] , 
        \b4_nUAi[893] , \b4_nUAi[894] , \b4_nUAi[895] , \b4_nUAi[896] , 
        \b4_nUAi[897] , \b4_nUAi[898] , \b4_nUAi[899] , \b4_nUAi[900] , 
        \b4_nUAi[901] , \b4_nUAi[902] , \b4_nUAi[903] , \b4_nUAi[904] , 
        \b4_nUAi[905] , \b4_nUAi[906] , \b4_nUAi[907] , \b4_nUAi[908] , 
        \b4_nUAi[909] , \b4_nUAi[910] , \b4_nUAi[911] , \b4_nUAi[912] , 
        \b4_nUAi[913] , \b4_nUAi[914] , \b4_nUAi[915] , \b4_nUAi[916] , 
        \b4_nUAi[917] , \b4_nUAi[918] , \b4_nUAi[919] , \b4_nUAi[920] , 
        \b4_nUAi[921] , \b4_nUAi[922] , \b4_nUAi[923] , \b4_nUAi[924] , 
        \b4_nUAi[925] , \b4_nUAi[926] , \b4_nUAi[927] , \b4_nUAi[928] , 
        \b4_nUAi[929] , \b4_nUAi[930] , \b4_nUAi[931] , \b4_nUAi[932] , 
        \b4_nUAi[933] , \b4_nUAi[934] , \b4_nUAi[935] , \b4_nUAi[936] , 
        \b4_nUAi[937] , \b4_nUAi[938] , \b4_nUAi[939] , \b4_nUAi[940] , 
        \b4_nUAi[941] , \b4_nUAi[942] , \b4_nUAi[943] , \b4_nUAi[944] , 
        \b4_nUAi[945] , \b4_nUAi[946] , \b4_nUAi[947] , \b4_nUAi[948] , 
        \b4_nUAi[949] , \b4_nUAi[950] , \b4_nUAi[951] , \b4_nUAi[952] , 
        \b4_nUAi[953] , \b4_nUAi[954] , \b4_nUAi[955] , \b4_nUAi[956] , 
        \b4_nUAi[957] , \b4_nUAi[958] , \b4_nUAi[959] , \b4_nUAi[960] , 
        \b4_nUAi[961] , \b4_nUAi[962] , \b4_nUAi[963] , \b4_nUAi[964] , 
        \b4_nUAi[965] , \b4_nUAi[966] , \b4_nUAi[967] , \b4_nUAi[968] , 
        \b4_nUAi[969] , \b4_nUAi[970] , \b4_nUAi[971] , \b4_nUAi[972] , 
        \b4_nUAi[973] , \b4_nUAi[974] , \b4_nUAi[975] , \b4_nUAi[976] , 
        \b4_nUAi[977] , \b4_nUAi[978] , \b4_nUAi[979] , \b4_nUAi[980] , 
        \b4_nUAi[981] , \b4_nUAi[982] , \b4_nUAi[983] , \b4_nUAi[984] , 
        \b4_nUAi[985] , \b4_nUAi[986] , \b4_nUAi[987] , \b4_nUAi[988] , 
        \b4_nUAi[989] , \b4_nUAi[990] , \b4_nUAi[991] , \b4_nUAi[992] , 
        \b4_nUAi[993] , \b4_nUAi[994] , \b4_nUAi[995] , \b4_nUAi[996] , 
        \b4_nUAi[997] , \b4_nUAi[998] , \b4_nUAi[999] , 
        \b4_nUAi[1000] , \b4_nUAi[1001] , \b4_nUAi[1002] , 
        \b4_nUAi[1003] , \b4_nUAi[1004] , \b4_nUAi[1005] , 
        \b4_nUAi[1006] , \b4_nUAi[1007] , \b4_nUAi[1008] , 
        \b4_nUAi[1009] , \b4_nUAi[1010] , \b4_nUAi[1011] , 
        \b4_nUAi[1012] , \b4_nUAi[1013] , \b4_nUAi[1014] , 
        \b4_nUAi[1015] , \b4_nUAi[1016] , \b4_nUAi[1017] , 
        \b4_nUAi[1018] , \b4_nUAi[1019] , \b4_nUAi[1020] , 
        \b4_nUAi[1021] , \b4_nUAi[1022] , \b4_nUAi[1023] , 
        \b4_nUAi[1024] , \b4_nUAi[1025] , \b4_nUAi[1026] , 
        \b4_nUAi[1027] , \b4_nUAi[1028] , \b4_nUAi[1029] , 
        \b4_nUAi[1030] , \b4_nUAi[1031] , \b4_nUAi[1032] , 
        \b4_nUAi[1033] , \b4_nUAi[1034] , \b4_nUAi[1035] , 
        \b4_nUAi[1036] , \b4_nUAi[1037] , \b4_nUAi[1038] , 
        \b4_nUAi[1039] , \b4_nUAi[1040] , \b4_nUAi[1041] , 
        \b4_nUAi[1042] , \b4_nUAi[1043] , \b4_nUAi[1044] , 
        \b4_nUAi[1045] , \b4_nUAi[1046] , \b4_nUAi[1047] , 
        \b4_nUAi[1048] , \b4_nUAi[1049] , \b4_nUAi[1050] , 
        \b4_nUAi[1051] , \b4_nUAi[1052] , \b4_nUAi[1053] , 
        \b4_nUAi[1054] , \b4_nUAi[1055] , \b4_nUAi[1056] , 
        \b4_nUAi[1057] , \b4_nUAi[1058] , \b4_nUAi[1059] , 
        \b4_nUAi[1060] , \b4_nUAi[1061] , \b4_nUAi[1062] , 
        \b4_nUAi[1063] , \b4_nUAi[1064] , \b4_nUAi[1065] , 
        \b4_nUAi[1066] , \b4_nUAi[1067] , \b4_nUAi[1068] , 
        \b4_nUAi[1069] , \b4_nUAi[1070] , \b4_nUAi[1071] , 
        \b4_nUAi[1072] , \b4_nUAi[1073] , \b4_nUAi[1074] , 
        \b4_nUAi[1075] , \b4_nUAi[1076] , \b4_nUAi[1077] , 
        \b4_nUAi[1078] , \b4_nUAi[1079] , \b4_nUAi[1080] , 
        \b4_nUAi[1081] , \b4_nUAi[1082] , \b4_nUAi[1083] , 
        \b4_nUAi[1084] , \b4_nUAi[1085] , \b4_nUAi[1086] , 
        \b4_nUAi[1087] , \b4_nUAi[1088] , \b4_nUAi[1089] , 
        \b4_nUAi[1090] , \b4_nUAi[1091] , \b4_nUAi[1092] , 
        \b4_nUAi[1093] , \b4_nUAi[1094] , \b4_nUAi[1095] , 
        \b4_nUAi[1096] , \b4_nUAi[1097] , \b4_nUAi[1098] , 
        \b4_nUAi[1099] , \b4_nUAi[1100] , \b4_nUAi[1101] , 
        \b4_nUAi[1102] , \b4_nUAi[1103] , \b4_nUAi[1104] , 
        \b4_nUAi[1105] , \b4_nUAi[1106] , \b4_nUAi[1107] , 
        \b4_nUAi[1108] , \b4_nUAi[1109] , \b4_nUAi[1110] , 
        \b4_nUAi[1111] , \b4_nUAi[1112] , \b4_nUAi[1113] , 
        \b4_nUAi[1114] , \b4_nUAi[1115] , \b4_nUAi[1116] , 
        \b4_nUAi[1117] , \b4_nUAi[1118] , \b4_nUAi[1119] , 
        \b4_nUAi[1120] , \b4_nUAi[1121] , \b4_nUAi[1122] , 
        \b4_nUAi[1123] , \b4_nUAi[1124] , \b4_nUAi[1125] , 
        \b4_nUAi[1126] , \b4_nUAi[1127] , \b4_nUAi[1128] , 
        \b4_nUAi[1129] ;
    
    b5_nvmFL_1131s_x b5_PbrtL (.b4_nUAi({\b4_nUAi[1129] , 
        \b4_nUAi[1128] , \b4_nUAi[1127] , \b4_nUAi[1126] , 
        \b4_nUAi[1125] , \b4_nUAi[1124] , \b4_nUAi[1123] , 
        \b4_nUAi[1122] , \b4_nUAi[1121] , \b4_nUAi[1120] , 
        \b4_nUAi[1119] , \b4_nUAi[1118] , \b4_nUAi[1117] , 
        \b4_nUAi[1116] , \b4_nUAi[1115] , \b4_nUAi[1114] , 
        \b4_nUAi[1113] , \b4_nUAi[1112] , \b4_nUAi[1111] , 
        \b4_nUAi[1110] , \b4_nUAi[1109] , \b4_nUAi[1108] , 
        \b4_nUAi[1107] , \b4_nUAi[1106] , \b4_nUAi[1105] , 
        \b4_nUAi[1104] , \b4_nUAi[1103] , \b4_nUAi[1102] , 
        \b4_nUAi[1101] , \b4_nUAi[1100] , \b4_nUAi[1099] , 
        \b4_nUAi[1098] , \b4_nUAi[1097] , \b4_nUAi[1096] , 
        \b4_nUAi[1095] , \b4_nUAi[1094] , \b4_nUAi[1093] , 
        \b4_nUAi[1092] , \b4_nUAi[1091] , \b4_nUAi[1090] , 
        \b4_nUAi[1089] , \b4_nUAi[1088] , \b4_nUAi[1087] , 
        \b4_nUAi[1086] , \b4_nUAi[1085] , \b4_nUAi[1084] , 
        \b4_nUAi[1083] , \b4_nUAi[1082] , \b4_nUAi[1081] , 
        \b4_nUAi[1080] , \b4_nUAi[1079] , \b4_nUAi[1078] , 
        \b4_nUAi[1077] , \b4_nUAi[1076] , \b4_nUAi[1075] , 
        \b4_nUAi[1074] , \b4_nUAi[1073] , \b4_nUAi[1072] , 
        \b4_nUAi[1071] , \b4_nUAi[1070] , \b4_nUAi[1069] , 
        \b4_nUAi[1068] , \b4_nUAi[1067] , \b4_nUAi[1066] , 
        \b4_nUAi[1065] , \b4_nUAi[1064] , \b4_nUAi[1063] , 
        \b4_nUAi[1062] , \b4_nUAi[1061] , \b4_nUAi[1060] , 
        \b4_nUAi[1059] , \b4_nUAi[1058] , \b4_nUAi[1057] , 
        \b4_nUAi[1056] , \b4_nUAi[1055] , \b4_nUAi[1054] , 
        \b4_nUAi[1053] , \b4_nUAi[1052] , \b4_nUAi[1051] , 
        \b4_nUAi[1050] , \b4_nUAi[1049] , \b4_nUAi[1048] , 
        \b4_nUAi[1047] , \b4_nUAi[1046] , \b4_nUAi[1045] , 
        \b4_nUAi[1044] , \b4_nUAi[1043] , \b4_nUAi[1042] , 
        \b4_nUAi[1041] , \b4_nUAi[1040] , \b4_nUAi[1039] , 
        \b4_nUAi[1038] , \b4_nUAi[1037] , \b4_nUAi[1036] , 
        \b4_nUAi[1035] , \b4_nUAi[1034] , \b4_nUAi[1033] , 
        \b4_nUAi[1032] , \b4_nUAi[1031] , \b4_nUAi[1030] , 
        \b4_nUAi[1029] , \b4_nUAi[1028] , \b4_nUAi[1027] , 
        \b4_nUAi[1026] , \b4_nUAi[1025] , \b4_nUAi[1024] , 
        \b4_nUAi[1023] , \b4_nUAi[1022] , \b4_nUAi[1021] , 
        \b4_nUAi[1020] , \b4_nUAi[1019] , \b4_nUAi[1018] , 
        \b4_nUAi[1017] , \b4_nUAi[1016] , \b4_nUAi[1015] , 
        \b4_nUAi[1014] , \b4_nUAi[1013] , \b4_nUAi[1012] , 
        \b4_nUAi[1011] , \b4_nUAi[1010] , \b4_nUAi[1009] , 
        \b4_nUAi[1008] , \b4_nUAi[1007] , \b4_nUAi[1006] , 
        \b4_nUAi[1005] , \b4_nUAi[1004] , \b4_nUAi[1003] , 
        \b4_nUAi[1002] , \b4_nUAi[1001] , \b4_nUAi[1000] , 
        \b4_nUAi[999] , \b4_nUAi[998] , \b4_nUAi[997] , \b4_nUAi[996] , 
        \b4_nUAi[995] , \b4_nUAi[994] , \b4_nUAi[993] , \b4_nUAi[992] , 
        \b4_nUAi[991] , \b4_nUAi[990] , \b4_nUAi[989] , \b4_nUAi[988] , 
        \b4_nUAi[987] , \b4_nUAi[986] , \b4_nUAi[985] , \b4_nUAi[984] , 
        \b4_nUAi[983] , \b4_nUAi[982] , \b4_nUAi[981] , \b4_nUAi[980] , 
        \b4_nUAi[979] , \b4_nUAi[978] , \b4_nUAi[977] , \b4_nUAi[976] , 
        \b4_nUAi[975] , \b4_nUAi[974] , \b4_nUAi[973] , \b4_nUAi[972] , 
        \b4_nUAi[971] , \b4_nUAi[970] , \b4_nUAi[969] , \b4_nUAi[968] , 
        \b4_nUAi[967] , \b4_nUAi[966] , \b4_nUAi[965] , \b4_nUAi[964] , 
        \b4_nUAi[963] , \b4_nUAi[962] , \b4_nUAi[961] , \b4_nUAi[960] , 
        \b4_nUAi[959] , \b4_nUAi[958] , \b4_nUAi[957] , \b4_nUAi[956] , 
        \b4_nUAi[955] , \b4_nUAi[954] , \b4_nUAi[953] , \b4_nUAi[952] , 
        \b4_nUAi[951] , \b4_nUAi[950] , \b4_nUAi[949] , \b4_nUAi[948] , 
        \b4_nUAi[947] , \b4_nUAi[946] , \b4_nUAi[945] , \b4_nUAi[944] , 
        \b4_nUAi[943] , \b4_nUAi[942] , \b4_nUAi[941] , \b4_nUAi[940] , 
        \b4_nUAi[939] , \b4_nUAi[938] , \b4_nUAi[937] , \b4_nUAi[936] , 
        \b4_nUAi[935] , \b4_nUAi[934] , \b4_nUAi[933] , \b4_nUAi[932] , 
        \b4_nUAi[931] , \b4_nUAi[930] , \b4_nUAi[929] , \b4_nUAi[928] , 
        \b4_nUAi[927] , \b4_nUAi[926] , \b4_nUAi[925] , \b4_nUAi[924] , 
        \b4_nUAi[923] , \b4_nUAi[922] , \b4_nUAi[921] , \b4_nUAi[920] , 
        \b4_nUAi[919] , \b4_nUAi[918] , \b4_nUAi[917] , \b4_nUAi[916] , 
        \b4_nUAi[915] , \b4_nUAi[914] , \b4_nUAi[913] , \b4_nUAi[912] , 
        \b4_nUAi[911] , \b4_nUAi[910] , \b4_nUAi[909] , \b4_nUAi[908] , 
        \b4_nUAi[907] , \b4_nUAi[906] , \b4_nUAi[905] , \b4_nUAi[904] , 
        \b4_nUAi[903] , \b4_nUAi[902] , \b4_nUAi[901] , \b4_nUAi[900] , 
        \b4_nUAi[899] , \b4_nUAi[898] , \b4_nUAi[897] , \b4_nUAi[896] , 
        \b4_nUAi[895] , \b4_nUAi[894] , \b4_nUAi[893] , \b4_nUAi[892] , 
        \b4_nUAi[891] , \b4_nUAi[890] , \b4_nUAi[889] , \b4_nUAi[888] , 
        \b4_nUAi[887] , \b4_nUAi[886] , \b4_nUAi[885] , \b4_nUAi[884] , 
        \b4_nUAi[883] , \b4_nUAi[882] , \b4_nUAi[881] , \b4_nUAi[880] , 
        \b4_nUAi[879] , \b4_nUAi[878] , \b4_nUAi[877] , \b4_nUAi[876] , 
        \b4_nUAi[875] , \b4_nUAi[874] , \b4_nUAi[873] , \b4_nUAi[872] , 
        \b4_nUAi[871] , \b4_nUAi[870] , \b4_nUAi[869] , \b4_nUAi[868] , 
        \b4_nUAi[867] , \b4_nUAi[866] , \b4_nUAi[865] , \b4_nUAi[864] , 
        \b4_nUAi[863] , \b4_nUAi[862] , \b4_nUAi[861] , \b4_nUAi[860] , 
        \b4_nUAi[859] , \b4_nUAi[858] , \b4_nUAi[857] , \b4_nUAi[856] , 
        \b4_nUAi[855] , \b4_nUAi[854] , \b4_nUAi[853] , \b4_nUAi[852] , 
        \b4_nUAi[851] , \b4_nUAi[850] , \b4_nUAi[849] , \b4_nUAi[848] , 
        \b4_nUAi[847] , \b4_nUAi[846] , \b4_nUAi[845] , \b4_nUAi[844] , 
        \b4_nUAi[843] , \b4_nUAi[842] , \b4_nUAi[841] , \b4_nUAi[840] , 
        \b4_nUAi[839] , \b4_nUAi[838] , \b4_nUAi[837] , \b4_nUAi[836] , 
        \b4_nUAi[835] , \b4_nUAi[834] , \b4_nUAi[833] , \b4_nUAi[832] , 
        \b4_nUAi[831] , \b4_nUAi[830] , \b4_nUAi[829] , \b4_nUAi[828] , 
        \b4_nUAi[827] , \b4_nUAi[826] , \b4_nUAi[825] , \b4_nUAi[824] , 
        \b4_nUAi[823] , \b4_nUAi[822] , \b4_nUAi[821] , \b4_nUAi[820] , 
        \b4_nUAi[819] , \b4_nUAi[818] , \b4_nUAi[817] , \b4_nUAi[816] , 
        \b4_nUAi[815] , \b4_nUAi[814] , \b4_nUAi[813] , \b4_nUAi[812] , 
        \b4_nUAi[811] , \b4_nUAi[810] , \b4_nUAi[809] , \b4_nUAi[808] , 
        \b4_nUAi[807] , \b4_nUAi[806] , \b4_nUAi[805] , \b4_nUAi[804] , 
        \b4_nUAi[803] , \b4_nUAi[802] , \b4_nUAi[801] , \b4_nUAi[800] , 
        \b4_nUAi[799] , \b4_nUAi[798] , \b4_nUAi[797] , \b4_nUAi[796] , 
        \b4_nUAi[795] , \b4_nUAi[794] , \b4_nUAi[793] , \b4_nUAi[792] , 
        \b4_nUAi[791] , \b4_nUAi[790] , \b4_nUAi[789] , \b4_nUAi[788] , 
        \b4_nUAi[787] , \b4_nUAi[786] , \b4_nUAi[785] , \b4_nUAi[784] , 
        \b4_nUAi[783] , \b4_nUAi[782] , \b4_nUAi[781] , \b4_nUAi[780] , 
        \b4_nUAi[779] , \b4_nUAi[778] , \b4_nUAi[777] , \b4_nUAi[776] , 
        \b4_nUAi[775] , \b4_nUAi[774] , \b4_nUAi[773] , \b4_nUAi[772] , 
        \b4_nUAi[771] , \b4_nUAi[770] , \b4_nUAi[769] , \b4_nUAi[768] , 
        \b4_nUAi[767] , \b4_nUAi[766] , \b4_nUAi[765] , \b4_nUAi[764] , 
        \b4_nUAi[763] , \b4_nUAi[762] , \b4_nUAi[761] , \b4_nUAi[760] , 
        \b4_nUAi[759] , \b4_nUAi[758] , \b4_nUAi[757] , \b4_nUAi[756] , 
        \b4_nUAi[755] , \b4_nUAi[754] , \b4_nUAi[753] , \b4_nUAi[752] , 
        \b4_nUAi[751] , \b4_nUAi[750] , \b4_nUAi[749] , \b4_nUAi[748] , 
        \b4_nUAi[747] , \b4_nUAi[746] , \b4_nUAi[745] , \b4_nUAi[744] , 
        \b4_nUAi[743] , \b4_nUAi[742] , \b4_nUAi[741] , \b4_nUAi[740] , 
        \b4_nUAi[739] , \b4_nUAi[738] , \b4_nUAi[737] , \b4_nUAi[736] , 
        \b4_nUAi[735] , \b4_nUAi[734] , \b4_nUAi[733] , \b4_nUAi[732] , 
        \b4_nUAi[731] , \b4_nUAi[730] , \b4_nUAi[729] , \b4_nUAi[728] , 
        \b4_nUAi[727] , \b4_nUAi[726] , \b4_nUAi[725] , \b4_nUAi[724] , 
        \b4_nUAi[723] , \b4_nUAi[722] , \b4_nUAi[721] , \b4_nUAi[720] , 
        \b4_nUAi[719] , \b4_nUAi[718] , \b4_nUAi[717] , \b4_nUAi[716] , 
        \b4_nUAi[715] , \b4_nUAi[714] , \b4_nUAi[713] , \b4_nUAi[712] , 
        \b4_nUAi[711] , \b4_nUAi[710] , \b4_nUAi[709] , \b4_nUAi[708] , 
        \b4_nUAi[707] , \b4_nUAi[706] , \b4_nUAi[705] , \b4_nUAi[704] , 
        \b4_nUAi[703] , \b4_nUAi[702] , \b4_nUAi[701] , \b4_nUAi[700] , 
        \b4_nUAi[699] , \b4_nUAi[698] , \b4_nUAi[697] , \b4_nUAi[696] , 
        \b4_nUAi[695] , \b4_nUAi[694] , \b4_nUAi[693] , \b4_nUAi[692] , 
        \b4_nUAi[691] , \b4_nUAi[690] , \b4_nUAi[689] , \b4_nUAi[688] , 
        \b4_nUAi[687] , \b4_nUAi[686] , \b4_nUAi[685] , \b4_nUAi[684] , 
        \b4_nUAi[683] , \b4_nUAi[682] , \b4_nUAi[681] , \b4_nUAi[680] , 
        \b4_nUAi[679] , \b4_nUAi[678] , \b4_nUAi[677] , \b4_nUAi[676] , 
        \b4_nUAi[675] , \b4_nUAi[674] , \b4_nUAi[673] , \b4_nUAi[672] , 
        \b4_nUAi[671] , \b4_nUAi[670] , \b4_nUAi[669] , \b4_nUAi[668] , 
        \b4_nUAi[667] , \b4_nUAi[666] , \b4_nUAi[665] , \b4_nUAi[664] , 
        \b4_nUAi[663] , \b4_nUAi[662] , \b4_nUAi[661] , \b4_nUAi[660] , 
        \b4_nUAi[659] , \b4_nUAi[658] , \b4_nUAi[657] , \b4_nUAi[656] , 
        \b4_nUAi[655] , \b4_nUAi[654] , \b4_nUAi[653] , \b4_nUAi[652] , 
        \b4_nUAi[651] , \b4_nUAi[650] , \b4_nUAi[649] , \b4_nUAi[648] , 
        \b4_nUAi[647] , \b4_nUAi[646] , \b4_nUAi[645] , \b4_nUAi[644] , 
        \b4_nUAi[643] , \b4_nUAi[642] , \b4_nUAi[641] , \b4_nUAi[640] , 
        \b4_nUAi[639] , \b4_nUAi[638] , \b4_nUAi[637] , \b4_nUAi[636] , 
        \b4_nUAi[635] , \b4_nUAi[634] , \b4_nUAi[633] , \b4_nUAi[632] , 
        \b4_nUAi[631] , \b4_nUAi[630] , \b4_nUAi[629] , \b4_nUAi[628] , 
        \b4_nUAi[627] , \b4_nUAi[626] , \b4_nUAi[625] , \b4_nUAi[624] , 
        \b4_nUAi[623] , \b4_nUAi[622] , \b4_nUAi[621] , \b4_nUAi[620] , 
        \b4_nUAi[619] , \b4_nUAi[618] , \b4_nUAi[617] , \b4_nUAi[616] , 
        \b4_nUAi[615] , \b4_nUAi[614] , \b4_nUAi[613] , \b4_nUAi[612] , 
        \b4_nUAi[611] , \b4_nUAi[610] , \b4_nUAi[609] , \b4_nUAi[608] , 
        \b4_nUAi[607] , \b4_nUAi[606] , \b4_nUAi[605] , \b4_nUAi[604] , 
        \b4_nUAi[603] , \b4_nUAi[602] , \b4_nUAi[601] , \b4_nUAi[600] , 
        \b4_nUAi[599] , \b4_nUAi[598] , \b4_nUAi[597] , \b4_nUAi[596] , 
        \b4_nUAi[595] , \b4_nUAi[594] , \b4_nUAi[593] , \b4_nUAi[592] , 
        \b4_nUAi[591] , \b4_nUAi[590] , \b4_nUAi[589] , \b4_nUAi[588] , 
        \b4_nUAi[587] , \b4_nUAi[586] , \b4_nUAi[585] , \b4_nUAi[584] , 
        \b4_nUAi[583] , \b4_nUAi[582] , \b4_nUAi[581] , \b4_nUAi[580] , 
        \b4_nUAi[579] , \b4_nUAi[578] , \b4_nUAi[577] , \b4_nUAi[576] , 
        \b4_nUAi[575] , \b4_nUAi[574] , \b4_nUAi[573] , \b4_nUAi[572] , 
        \b4_nUAi[571] , \b4_nUAi[570] , \b4_nUAi[569] , \b4_nUAi[568] , 
        \b4_nUAi[567] , \b4_nUAi[566] , \b4_nUAi[565] , \b4_nUAi[564] , 
        \b4_nUAi[563] , \b4_nUAi[562] , \b4_nUAi[561] , \b4_nUAi[560] , 
        \b4_nUAi[559] , \b4_nUAi[558] , \b4_nUAi[557] , \b4_nUAi[556] , 
        \b4_nUAi[555] , \b4_nUAi[554] , \b4_nUAi[553] , \b4_nUAi[552] , 
        \b4_nUAi[551] , \b4_nUAi[550] , \b4_nUAi[549] , \b4_nUAi[548] , 
        \b4_nUAi[547] , \b4_nUAi[546] , \b4_nUAi[545] , \b4_nUAi[544] , 
        \b4_nUAi[543] , \b4_nUAi[542] , \b4_nUAi[541] , \b4_nUAi[540] , 
        \b4_nUAi[539] , \b4_nUAi[538] , \b4_nUAi[537] , \b4_nUAi[536] , 
        \b4_nUAi[535] , \b4_nUAi[534] , \b4_nUAi[533] , \b4_nUAi[532] , 
        \b4_nUAi[531] , \b4_nUAi[530] , \b4_nUAi[529] , \b4_nUAi[528] , 
        \b4_nUAi[527] , \b4_nUAi[526] , \b4_nUAi[525] , \b4_nUAi[524] , 
        \b4_nUAi[523] , \b4_nUAi[522] , \b4_nUAi[521] , \b4_nUAi[520] , 
        \b4_nUAi[519] , \b4_nUAi[518] , \b4_nUAi[517] , \b4_nUAi[516] , 
        \b4_nUAi[515] , \b4_nUAi[514] , \b4_nUAi[513] , \b4_nUAi[512] , 
        \b4_nUAi[511] , \b4_nUAi[510] , \b4_nUAi[509] , \b4_nUAi[508] , 
        \b4_nUAi[507] , \b4_nUAi[506] , \b4_nUAi[505] , \b4_nUAi[504] , 
        \b4_nUAi[503] , \b4_nUAi[502] , \b4_nUAi[501] , \b4_nUAi[500] , 
        \b4_nUAi[499] , \b4_nUAi[498] , \b4_nUAi[497] , \b4_nUAi[496] , 
        \b4_nUAi[495] , \b4_nUAi[494] , \b4_nUAi[493] , \b4_nUAi[492] , 
        \b4_nUAi[491] , \b4_nUAi[490] , \b4_nUAi[489] , \b4_nUAi[488] , 
        \b4_nUAi[487] , \b4_nUAi[486] , \b4_nUAi[485] , \b4_nUAi[484] , 
        \b4_nUAi[483] , \b4_nUAi[482] , \b4_nUAi[481] , \b4_nUAi[480] , 
        \b4_nUAi[479] , \b4_nUAi[478] , \b4_nUAi[477] , \b4_nUAi[476] , 
        \b4_nUAi[475] , \b4_nUAi[474] , \b4_nUAi[473] , \b4_nUAi[472] , 
        \b4_nUAi[471] , \b4_nUAi[470] , \b4_nUAi[469] , \b4_nUAi[468] , 
        \b4_nUAi[467] , \b4_nUAi[466] , \b4_nUAi[465] , \b4_nUAi[464] , 
        \b4_nUAi[463] , \b4_nUAi[462] , \b4_nUAi[461] , \b4_nUAi[460] , 
        \b4_nUAi[459] , \b4_nUAi[458] , \b4_nUAi[457] , \b4_nUAi[456] , 
        \b4_nUAi[455] , \b4_nUAi[454] , \b4_nUAi[453] , \b4_nUAi[452] , 
        \b4_nUAi[451] , \b4_nUAi[450] , \b4_nUAi[449] , \b4_nUAi[448] , 
        \b4_nUAi[447] , \b4_nUAi[446] , \b4_nUAi[445] , \b4_nUAi[444] , 
        \b4_nUAi[443] , \b4_nUAi[442] , \b4_nUAi[441] , \b4_nUAi[440] , 
        \b4_nUAi[439] , \b4_nUAi[438] , \b4_nUAi[437] , \b4_nUAi[436] , 
        \b4_nUAi[435] , \b4_nUAi[434] , \b4_nUAi[433] , \b4_nUAi[432] , 
        \b4_nUAi[431] , \b4_nUAi[430] , \b4_nUAi[429] , \b4_nUAi[428] , 
        \b4_nUAi[427] , \b4_nUAi[426] , \b4_nUAi[425] , \b4_nUAi[424] , 
        \b4_nUAi[423] , \b4_nUAi[422] , \b4_nUAi[421] , \b4_nUAi[420] , 
        \b4_nUAi[419] , \b4_nUAi[418] , \b4_nUAi[417] , \b4_nUAi[416] , 
        \b4_nUAi[415] , \b4_nUAi[414] , \b4_nUAi[413] , \b4_nUAi[412] , 
        \b4_nUAi[411] , \b4_nUAi[410] , \b4_nUAi[409] , \b4_nUAi[408] , 
        \b4_nUAi[407] , \b4_nUAi[406] , \b4_nUAi[405] , \b4_nUAi[404] , 
        \b4_nUAi[403] , \b4_nUAi[402] , \b4_nUAi[401] , \b4_nUAi[400] , 
        \b4_nUAi[399] , \b4_nUAi[398] , \b4_nUAi[397] , \b4_nUAi[396] , 
        \b4_nUAi[395] , \b4_nUAi[394] , \b4_nUAi[393] , \b4_nUAi[392] , 
        \b4_nUAi[391] , \b4_nUAi[390] , \b4_nUAi[389] , \b4_nUAi[388] , 
        \b4_nUAi[387] , \b4_nUAi[386] , \b4_nUAi[385] , \b4_nUAi[384] , 
        \b4_nUAi[383] , \b4_nUAi[382] , \b4_nUAi[381] , \b4_nUAi[380] , 
        \b4_nUAi[379] , \b4_nUAi[378] , \b4_nUAi[377] , \b4_nUAi[376] , 
        \b4_nUAi[375] , \b4_nUAi[374] , \b4_nUAi[373] , \b4_nUAi[372] , 
        \b4_nUAi[371] , \b4_nUAi[370] , \b4_nUAi[369] , \b4_nUAi[368] , 
        \b4_nUAi[367] , \b4_nUAi[366] , \b4_nUAi[365] , \b4_nUAi[364] , 
        \b4_nUAi[363] , \b4_nUAi[362] , \b4_nUAi[361] , \b4_nUAi[360] , 
        \b4_nUAi[359] , \b4_nUAi[358] , \b4_nUAi[357] , \b4_nUAi[356] , 
        \b4_nUAi[355] , \b4_nUAi[354] , \b4_nUAi[353] , \b4_nUAi[352] , 
        \b4_nUAi[351] , \b4_nUAi[350] , \b4_nUAi[349] , \b4_nUAi[348] , 
        \b4_nUAi[347] , \b4_nUAi[346] , \b4_nUAi[345] , \b4_nUAi[344] , 
        \b4_nUAi[343] , \b4_nUAi[342] , \b4_nUAi[341] , \b4_nUAi[340] , 
        \b4_nUAi[339] , \b4_nUAi[338] , \b4_nUAi[337] , \b4_nUAi[336] , 
        \b4_nUAi[335] , \b4_nUAi[334] , \b4_nUAi[333] , \b4_nUAi[332] , 
        \b4_nUAi[331] , \b4_nUAi[330] , \b4_nUAi[329] , \b4_nUAi[328] , 
        \b4_nUAi[327] , \b4_nUAi[326] , \b4_nUAi[325] , \b4_nUAi[324] , 
        \b4_nUAi[323] , \b4_nUAi[322] , \b4_nUAi[321] , \b4_nUAi[320] , 
        \b4_nUAi[319] , \b4_nUAi[318] , \b4_nUAi[317] , \b4_nUAi[316] , 
        \b4_nUAi[315] , \b4_nUAi[314] , \b4_nUAi[313] , \b4_nUAi[312] , 
        \b4_nUAi[311] , \b4_nUAi[310] , \b4_nUAi[309] , \b4_nUAi[308] , 
        \b4_nUAi[307] , \b4_nUAi[306] , \b4_nUAi[305] , \b4_nUAi[304] , 
        \b4_nUAi[303] , \b4_nUAi[302] , \b4_nUAi[301] , \b4_nUAi[300] , 
        \b4_nUAi[299] , \b4_nUAi[298] , \b4_nUAi[297] , \b4_nUAi[296] , 
        \b4_nUAi[295] , \b4_nUAi[294] , \b4_nUAi[293] , \b4_nUAi[292] , 
        \b4_nUAi[291] , \b4_nUAi[290] , \b4_nUAi[289] , \b4_nUAi[288] , 
        \b4_nUAi[287] , \b4_nUAi[286] , \b4_nUAi[285] , \b4_nUAi[284] , 
        \b4_nUAi[283] , \b4_nUAi[282] , \b4_nUAi[281] , \b4_nUAi[280] , 
        \b4_nUAi[279] , \b4_nUAi[278] , \b4_nUAi[277] , \b4_nUAi[276] , 
        \b4_nUAi[275] , \b4_nUAi[274] , \b4_nUAi[273] , \b4_nUAi[272] , 
        \b4_nUAi[271] , \b4_nUAi[270] , \b4_nUAi[269] , \b4_nUAi[268] , 
        \b4_nUAi[267] , \b4_nUAi[266] , \b4_nUAi[265] , \b4_nUAi[264] , 
        \b4_nUAi[263] , \b4_nUAi[262] , \b4_nUAi[261] , \b4_nUAi[260] , 
        \b4_nUAi[259] , \b4_nUAi[258] , \b4_nUAi[257] , \b4_nUAi[256] , 
        \b4_nUAi[255] , \b4_nUAi[254] , \b4_nUAi[253] , \b4_nUAi[252] , 
        \b4_nUAi[251] , \b4_nUAi[250] , \b4_nUAi[249] , \b4_nUAi[248] , 
        \b4_nUAi[247] , \b4_nUAi[246] , \b4_nUAi[245] , \b4_nUAi[244] , 
        \b4_nUAi[243] , \b4_nUAi[242] , \b4_nUAi[241] , \b4_nUAi[240] , 
        \b4_nUAi[239] , \b4_nUAi[238] , \b4_nUAi[237] , \b4_nUAi[236] , 
        \b4_nUAi[235] , \b4_nUAi[234] , \b4_nUAi[233] , \b4_nUAi[232] , 
        \b4_nUAi[231] , \b4_nUAi[230] , \b4_nUAi[229] , \b4_nUAi[228] , 
        \b4_nUAi[227] , \b4_nUAi[226] , \b4_nUAi[225] , \b4_nUAi[224] , 
        \b4_nUAi[223] , \b4_nUAi[222] , \b4_nUAi[221] , \b4_nUAi[220] , 
        \b4_nUAi[219] , \b4_nUAi[218] , \b4_nUAi[217] , \b4_nUAi[216] , 
        \b4_nUAi[215] , \b4_nUAi[214] , \b4_nUAi[213] , \b4_nUAi[212] , 
        \b4_nUAi[211] , \b4_nUAi[210] , \b4_nUAi[209] , \b4_nUAi[208] , 
        \b4_nUAi[207] , \b4_nUAi[206] , \b4_nUAi[205] , \b4_nUAi[204] , 
        \b4_nUAi[203] , \b4_nUAi[202] , \b4_nUAi[201] , \b4_nUAi[200] , 
        \b4_nUAi[199] , \b4_nUAi[198] , \b4_nUAi[197] , \b4_nUAi[196] , 
        \b4_nUAi[195] , \b4_nUAi[194] , \b4_nUAi[193] , \b4_nUAi[192] , 
        \b4_nUAi[191] , \b4_nUAi[190] , \b4_nUAi[189] , \b4_nUAi[188] , 
        \b4_nUAi[187] , \b4_nUAi[186] , \b4_nUAi[185] , \b4_nUAi[184] , 
        \b4_nUAi[183] , \b4_nUAi[182] , \b4_nUAi[181] , \b4_nUAi[180] , 
        \b4_nUAi[179] , \b4_nUAi[178] , \b4_nUAi[177] , \b4_nUAi[176] , 
        \b4_nUAi[175] , \b4_nUAi[174] , \b4_nUAi[173] , \b4_nUAi[172] , 
        \b4_nUAi[171] , \b4_nUAi[170] , \b4_nUAi[169] , \b4_nUAi[168] , 
        \b4_nUAi[167] , \b4_nUAi[166] , \b4_nUAi[165] , \b4_nUAi[164] , 
        \b4_nUAi[163] , \b4_nUAi[162] , \b4_nUAi[161] , \b4_nUAi[160] , 
        \b4_nUAi[159] , \b4_nUAi[158] , \b4_nUAi[157] , \b4_nUAi[156] , 
        \b4_nUAi[155] , \b4_nUAi[154] , \b4_nUAi[153] , \b4_nUAi[152] , 
        \b4_nUAi[151] , \b4_nUAi[150] , \b4_nUAi[149] , \b4_nUAi[148] , 
        \b4_nUAi[147] , \b4_nUAi[146] , \b4_nUAi[145] , \b4_nUAi[144] , 
        \b4_nUAi[143] , \b4_nUAi[142] , \b4_nUAi[141] , \b4_nUAi[140] , 
        \b4_nUAi[139] , \b4_nUAi[138] , \b4_nUAi[137] , \b4_nUAi[136] , 
        \b4_nUAi[135] , \b4_nUAi[134] , \b4_nUAi[133] , \b4_nUAi[132] , 
        \b4_nUAi[131] , \b4_nUAi[130] , \b4_nUAi[129] , \b4_nUAi[128] , 
        \b4_nUAi[127] , \b4_nUAi[126] , \b4_nUAi[125] , \b4_nUAi[124] , 
        \b4_nUAi[123] , \b4_nUAi[122] , \b4_nUAi[121] , \b4_nUAi[120] , 
        \b4_nUAi[119] , \b4_nUAi[118] , \b4_nUAi[117] , \b4_nUAi[116] , 
        \b4_nUAi[115] , \b4_nUAi[114] , \b4_nUAi[113] , \b4_nUAi[112] , 
        \b4_nUAi[111] , \b4_nUAi[110] , \b4_nUAi[109] , \b4_nUAi[108] , 
        \b4_nUAi[107] , \b4_nUAi[106] , \b4_nUAi[105] , \b4_nUAi[104] , 
        \b4_nUAi[103] , \b4_nUAi[102] , \b4_nUAi[101] , \b4_nUAi[100] , 
        \b4_nUAi[99] , \b4_nUAi[98] , \b4_nUAi[97] , \b4_nUAi[96] , 
        \b4_nUAi[95] , \b4_nUAi[94] , \b4_nUAi[93] , \b4_nUAi[92] , 
        \b4_nUAi[91] , \b4_nUAi[90] , \b4_nUAi[89] , \b4_nUAi[88] , 
        \b4_nUAi[87] , \b4_nUAi[86] , \b4_nUAi[85] , \b4_nUAi[84] , 
        \b4_nUAi[83] , \b4_nUAi[82] , \b4_nUAi[81] , \b4_nUAi[80] , 
        \b4_nUAi[79] , \b4_nUAi[78] , \b4_nUAi[77] , \b4_nUAi[76] , 
        \b4_nUAi[75] , \b4_nUAi[74] , \b4_nUAi[73] , \b4_nUAi[72] , 
        \b4_nUAi[71] , \b4_nUAi[70] , \b4_nUAi[69] , \b4_nUAi[68] , 
        \b4_nUAi[67] , \b4_nUAi[66] , \b4_nUAi[65] , \b4_nUAi[64] , 
        \b4_nUAi[63] , \b4_nUAi[62] , \b4_nUAi[61] , \b4_nUAi[60] , 
        \b4_nUAi[59] , \b4_nUAi[58] , \b4_nUAi[57] , \b4_nUAi[56] , 
        \b4_nUAi[55] , \b4_nUAi[54] , \b4_nUAi[53] , \b4_nUAi[52] , 
        \b4_nUAi[51] , \b4_nUAi[50] , \b4_nUAi[49] , \b4_nUAi[48] , 
        \b4_nUAi[47] , \b4_nUAi[46] , \b4_nUAi[45] , \b4_nUAi[44] , 
        \b4_nUAi[43] , \b4_nUAi[42] , \b4_nUAi[41] , \b4_nUAi[40] , 
        \b4_nUAi[39] , \b4_nUAi[38] , \b4_nUAi[37] , \b4_nUAi[36] , 
        \b4_nUAi[35] , \b4_nUAi[34] , \b4_nUAi[33] , \b4_nUAi[32] , 
        \b4_nUAi[31] , \b4_nUAi[30] , \b4_nUAi[29] , \b4_nUAi[28] , 
        \b4_nUAi[27] , \b4_nUAi[26] , \b4_nUAi[25] , \b4_nUAi[24] , 
        \b4_nUAi[23] , \b4_nUAi[22] , \b4_nUAi[21] , \b4_nUAi[20] , 
        \b4_nUAi[19] , \b4_nUAi[18] , \b4_nUAi[17] , \b4_nUAi[16] , 
        \b4_nUAi[15] , \b4_nUAi[14] , \b4_nUAi[13] , \b4_nUAi[12] , 
        \b4_nUAi[11] , \b4_nUAi[10] , \b4_nUAi[9] , \b4_nUAi[8] , 
        \b4_nUAi[7] , \b4_nUAi[6] , \b4_nUAi[5] , \b4_nUAi[4] , 
        \b4_nUAi[3] , \b4_nUAi[2] , \b4_nUAi[1] , \b4_nUAi[0] }), 
        .IICE_comm2iice({IICE_comm2iice[11], IICE_comm2iice[10]}), 
        .b4_PLyF(b4_PLyF), .b7_PSyi3wy(b7_PSyi3wy), .b8_PSyiBgYG(
        b8_PSyiBgYG));
    VCC VCC (.Y(VCC_net_1));
    b11_PSyil9s1fkT_x b7_PbTtl9G (.mdiclink_reg({mdiclink_reg[376], 
        mdiclink_reg[375], mdiclink_reg[374], mdiclink_reg[373], 
        mdiclink_reg[372], mdiclink_reg[371], mdiclink_reg[370], 
        mdiclink_reg[369], mdiclink_reg[368], mdiclink_reg[367], 
        mdiclink_reg[366], mdiclink_reg[365], mdiclink_reg[364], 
        mdiclink_reg[363], mdiclink_reg[362], mdiclink_reg[361], 
        mdiclink_reg[360], mdiclink_reg[359], mdiclink_reg[358], 
        mdiclink_reg[357], mdiclink_reg[356], mdiclink_reg[355], 
        mdiclink_reg[354], mdiclink_reg[353], mdiclink_reg[352], 
        mdiclink_reg[351], mdiclink_reg[350], mdiclink_reg[349], 
        mdiclink_reg[348], mdiclink_reg[347], mdiclink_reg[346], 
        mdiclink_reg[345], mdiclink_reg[344], mdiclink_reg[343], 
        mdiclink_reg[342], mdiclink_reg[341], mdiclink_reg[340], 
        mdiclink_reg[339], mdiclink_reg[338], mdiclink_reg[337], 
        mdiclink_reg[336], mdiclink_reg[335], mdiclink_reg[334], 
        mdiclink_reg[333], mdiclink_reg[332], mdiclink_reg[331], 
        mdiclink_reg[330], mdiclink_reg[329], mdiclink_reg[328], 
        mdiclink_reg[327], mdiclink_reg[326], mdiclink_reg[325], 
        mdiclink_reg[324], mdiclink_reg[323], mdiclink_reg[322], 
        mdiclink_reg[321], mdiclink_reg[320], mdiclink_reg[319], 
        mdiclink_reg[318], mdiclink_reg[317], mdiclink_reg[316], 
        mdiclink_reg[315], mdiclink_reg[314], mdiclink_reg[313], 
        mdiclink_reg[312], mdiclink_reg[311], mdiclink_reg[310], 
        mdiclink_reg[309], mdiclink_reg[308], mdiclink_reg[307], 
        mdiclink_reg[306], mdiclink_reg[305], mdiclink_reg[304], 
        mdiclink_reg[303], mdiclink_reg[302], mdiclink_reg[301], 
        mdiclink_reg[300], mdiclink_reg[299], mdiclink_reg[298], 
        mdiclink_reg[297], mdiclink_reg[296], mdiclink_reg[295], 
        mdiclink_reg[294], mdiclink_reg[293], mdiclink_reg[292], 
        mdiclink_reg[291], mdiclink_reg[290], mdiclink_reg[289], 
        mdiclink_reg[288], mdiclink_reg[287], mdiclink_reg[286], 
        mdiclink_reg[285], mdiclink_reg[284], mdiclink_reg[283], 
        mdiclink_reg[282], mdiclink_reg[281], mdiclink_reg[280], 
        mdiclink_reg[279], mdiclink_reg[278], mdiclink_reg[277], 
        mdiclink_reg[276], mdiclink_reg[275], mdiclink_reg[274], 
        mdiclink_reg[273], mdiclink_reg[272], mdiclink_reg[271], 
        mdiclink_reg[270], mdiclink_reg[269], mdiclink_reg[268], 
        mdiclink_reg[267], mdiclink_reg[266], mdiclink_reg[265], 
        mdiclink_reg[264], mdiclink_reg[263], mdiclink_reg[262], 
        mdiclink_reg[261], mdiclink_reg[260], mdiclink_reg[259], 
        mdiclink_reg[258], mdiclink_reg[257], mdiclink_reg[256], 
        mdiclink_reg[255], mdiclink_reg[254], mdiclink_reg[253], 
        mdiclink_reg[252], mdiclink_reg[251], mdiclink_reg[250], 
        mdiclink_reg[249], mdiclink_reg[248], mdiclink_reg[247], 
        mdiclink_reg[246], mdiclink_reg[245], mdiclink_reg[244], 
        mdiclink_reg[243], mdiclink_reg[242], mdiclink_reg[241], 
        mdiclink_reg[240], mdiclink_reg[239], mdiclink_reg[238], 
        mdiclink_reg[237], mdiclink_reg[236], mdiclink_reg[235], 
        mdiclink_reg[234], mdiclink_reg[233], mdiclink_reg[232], 
        mdiclink_reg[231], mdiclink_reg[230], mdiclink_reg[229], 
        mdiclink_reg[228], mdiclink_reg[227], mdiclink_reg[226], 
        mdiclink_reg[225], mdiclink_reg[224], mdiclink_reg[223], 
        mdiclink_reg[222], mdiclink_reg[221], mdiclink_reg[220], 
        mdiclink_reg[219], mdiclink_reg[218], mdiclink_reg[217], 
        mdiclink_reg[216], mdiclink_reg[215], mdiclink_reg[214], 
        mdiclink_reg[213], mdiclink_reg[212], mdiclink_reg[211], 
        mdiclink_reg[210], mdiclink_reg[209], mdiclink_reg[208], 
        mdiclink_reg[207], mdiclink_reg[206], mdiclink_reg[205], 
        mdiclink_reg[204], mdiclink_reg[203], mdiclink_reg[202], 
        mdiclink_reg[201], mdiclink_reg[200], mdiclink_reg[199], 
        mdiclink_reg[198], mdiclink_reg[197], mdiclink_reg[196], 
        mdiclink_reg[195], mdiclink_reg[194], mdiclink_reg[193], 
        mdiclink_reg[192], mdiclink_reg[191], mdiclink_reg[190], 
        mdiclink_reg[189], mdiclink_reg[188], mdiclink_reg[187], 
        mdiclink_reg[186], mdiclink_reg[185], mdiclink_reg[184], 
        mdiclink_reg[183], mdiclink_reg[182], mdiclink_reg[181], 
        mdiclink_reg[180], mdiclink_reg[179], mdiclink_reg[178], 
        mdiclink_reg[177], mdiclink_reg[176], mdiclink_reg[175], 
        mdiclink_reg[174], mdiclink_reg[173], mdiclink_reg[172], 
        mdiclink_reg[171], mdiclink_reg[170], mdiclink_reg[169], 
        mdiclink_reg[168], mdiclink_reg[167], mdiclink_reg[166], 
        mdiclink_reg[165], mdiclink_reg[164], mdiclink_reg[163], 
        mdiclink_reg[162], mdiclink_reg[161], mdiclink_reg[160], 
        mdiclink_reg[159], mdiclink_reg[158], mdiclink_reg[157], 
        mdiclink_reg[156], mdiclink_reg[155], mdiclink_reg[154], 
        mdiclink_reg[153], mdiclink_reg[152], mdiclink_reg[151], 
        mdiclink_reg[150], mdiclink_reg[149], mdiclink_reg[148], 
        mdiclink_reg[147], mdiclink_reg[146], mdiclink_reg[145], 
        mdiclink_reg[144], mdiclink_reg[143], mdiclink_reg[142], 
        mdiclink_reg[141], mdiclink_reg[140], mdiclink_reg[139], 
        mdiclink_reg[138], mdiclink_reg[137], mdiclink_reg[136], 
        mdiclink_reg[135], mdiclink_reg[134], mdiclink_reg[133], 
        mdiclink_reg[132], mdiclink_reg[131], mdiclink_reg[130], 
        mdiclink_reg[129], mdiclink_reg[128], mdiclink_reg[127], 
        mdiclink_reg[126], mdiclink_reg[125], mdiclink_reg[124], 
        mdiclink_reg[123], mdiclink_reg[122], mdiclink_reg[121], 
        mdiclink_reg[120], mdiclink_reg[119], mdiclink_reg[118], 
        mdiclink_reg[117], mdiclink_reg[116], mdiclink_reg[115], 
        mdiclink_reg[114], mdiclink_reg[113], mdiclink_reg[112], 
        mdiclink_reg[111], mdiclink_reg[110], mdiclink_reg[109], 
        mdiclink_reg[108], mdiclink_reg[107], mdiclink_reg[106], 
        mdiclink_reg[105], mdiclink_reg[104], mdiclink_reg[103], 
        mdiclink_reg[102], mdiclink_reg[101], mdiclink_reg[100], 
        mdiclink_reg[99], mdiclink_reg[98], mdiclink_reg[97], 
        mdiclink_reg[96], mdiclink_reg[95], mdiclink_reg[94], 
        mdiclink_reg[93], mdiclink_reg[92], mdiclink_reg[91], 
        mdiclink_reg[90], mdiclink_reg[89], mdiclink_reg[88], 
        mdiclink_reg[87], mdiclink_reg[86], mdiclink_reg[85], 
        mdiclink_reg[84], mdiclink_reg[83], mdiclink_reg[82], 
        mdiclink_reg[81], mdiclink_reg[80], mdiclink_reg[79], 
        mdiclink_reg[78], mdiclink_reg[77], mdiclink_reg[76], 
        mdiclink_reg[75], mdiclink_reg[74], mdiclink_reg[73], 
        mdiclink_reg[72], mdiclink_reg[71], mdiclink_reg[70], 
        mdiclink_reg[69], mdiclink_reg[68], mdiclink_reg[67], 
        mdiclink_reg[66], mdiclink_reg[65], mdiclink_reg[64], 
        mdiclink_reg[63], mdiclink_reg[62], mdiclink_reg[61], 
        mdiclink_reg[60], mdiclink_reg[59], mdiclink_reg[58], 
        mdiclink_reg[57], mdiclink_reg[56], mdiclink_reg[55], 
        mdiclink_reg[54], mdiclink_reg[53], mdiclink_reg[52], 
        mdiclink_reg[51], mdiclink_reg[50], mdiclink_reg[49], 
        mdiclink_reg[48], mdiclink_reg[47], mdiclink_reg[46], 
        mdiclink_reg[45], mdiclink_reg[44], mdiclink_reg[43], 
        mdiclink_reg[42], mdiclink_reg[41], mdiclink_reg[40], 
        mdiclink_reg[39], mdiclink_reg[38], mdiclink_reg[37], 
        mdiclink_reg[36], mdiclink_reg[35], mdiclink_reg[34], 
        mdiclink_reg[33], mdiclink_reg[32], mdiclink_reg[31], 
        mdiclink_reg[30], mdiclink_reg[29], mdiclink_reg[28], 
        mdiclink_reg[27], mdiclink_reg[26], mdiclink_reg[25], 
        mdiclink_reg[24], mdiclink_reg[23], mdiclink_reg[22], 
        mdiclink_reg[21], mdiclink_reg[20], mdiclink_reg[19], 
        mdiclink_reg[18], mdiclink_reg[17], mdiclink_reg[16], 
        mdiclink_reg[15], mdiclink_reg[14], mdiclink_reg[13], 
        mdiclink_reg[12], mdiclink_reg[11], mdiclink_reg[10], 
        mdiclink_reg[9], mdiclink_reg[8], mdiclink_reg[7], 
        mdiclink_reg[6], mdiclink_reg[5], mdiclink_reg[4], 
        mdiclink_reg[3], mdiclink_reg[2], mdiclink_reg[1], 
        mdiclink_reg[0]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[376], 
        b11_OFWNT9L_8tZ[375], b11_OFWNT9L_8tZ[374], 
        b11_OFWNT9L_8tZ[373], b11_OFWNT9L_8tZ[372], 
        b11_OFWNT9L_8tZ[371], b11_OFWNT9L_8tZ[370], 
        b11_OFWNT9L_8tZ[369], b11_OFWNT9L_8tZ[368], 
        b11_OFWNT9L_8tZ[367], b11_OFWNT9L_8tZ[366], 
        b11_OFWNT9L_8tZ[365], b11_OFWNT9L_8tZ[364], 
        b11_OFWNT9L_8tZ[363], b11_OFWNT9L_8tZ[362], 
        b11_OFWNT9L_8tZ[361], b11_OFWNT9L_8tZ[360], 
        b11_OFWNT9L_8tZ[359], b11_OFWNT9L_8tZ[358], 
        b11_OFWNT9L_8tZ[357], b11_OFWNT9L_8tZ[356], 
        b11_OFWNT9L_8tZ[355], b11_OFWNT9L_8tZ[354], 
        b11_OFWNT9L_8tZ[353], b11_OFWNT9L_8tZ[352], 
        b11_OFWNT9L_8tZ[351], b11_OFWNT9L_8tZ[350], 
        b11_OFWNT9L_8tZ[349], b11_OFWNT9L_8tZ[348], 
        b11_OFWNT9L_8tZ[347], b11_OFWNT9L_8tZ[346], 
        b11_OFWNT9L_8tZ[345], b11_OFWNT9L_8tZ[344], 
        b11_OFWNT9L_8tZ[343], b11_OFWNT9L_8tZ[342], 
        b11_OFWNT9L_8tZ[341], b11_OFWNT9L_8tZ[340], 
        b11_OFWNT9L_8tZ[339], b11_OFWNT9L_8tZ[338], 
        b11_OFWNT9L_8tZ[337], b11_OFWNT9L_8tZ[336], 
        b11_OFWNT9L_8tZ[335], b11_OFWNT9L_8tZ[334], 
        b11_OFWNT9L_8tZ[333], b11_OFWNT9L_8tZ[332], 
        b11_OFWNT9L_8tZ[331], b11_OFWNT9L_8tZ[330], 
        b11_OFWNT9L_8tZ[329], b11_OFWNT9L_8tZ[328], 
        b11_OFWNT9L_8tZ[327], b11_OFWNT9L_8tZ[326], 
        b11_OFWNT9L_8tZ[325], b11_OFWNT9L_8tZ[324], 
        b11_OFWNT9L_8tZ[323], b11_OFWNT9L_8tZ[322], 
        b11_OFWNT9L_8tZ[321], b11_OFWNT9L_8tZ[320], 
        b11_OFWNT9L_8tZ[319], b11_OFWNT9L_8tZ[318], 
        b11_OFWNT9L_8tZ[317], b11_OFWNT9L_8tZ[316], 
        b11_OFWNT9L_8tZ[315], b11_OFWNT9L_8tZ[314], 
        b11_OFWNT9L_8tZ[313], b11_OFWNT9L_8tZ[312], 
        b11_OFWNT9L_8tZ[311], b11_OFWNT9L_8tZ[310], 
        b11_OFWNT9L_8tZ[309], b11_OFWNT9L_8tZ[308], 
        b11_OFWNT9L_8tZ[307], b11_OFWNT9L_8tZ[306], 
        b11_OFWNT9L_8tZ[305], b11_OFWNT9L_8tZ[304], 
        b11_OFWNT9L_8tZ[303], b11_OFWNT9L_8tZ[302], 
        b11_OFWNT9L_8tZ[301], b11_OFWNT9L_8tZ[300], 
        b11_OFWNT9L_8tZ[299], b11_OFWNT9L_8tZ[298], 
        b11_OFWNT9L_8tZ[297], b11_OFWNT9L_8tZ[296], 
        b11_OFWNT9L_8tZ[295], b11_OFWNT9L_8tZ[294], 
        b11_OFWNT9L_8tZ[293], b11_OFWNT9L_8tZ[292], 
        b11_OFWNT9L_8tZ[291], b11_OFWNT9L_8tZ[290], 
        b11_OFWNT9L_8tZ[289], b11_OFWNT9L_8tZ[288], 
        b11_OFWNT9L_8tZ[287], b11_OFWNT9L_8tZ[286], 
        b11_OFWNT9L_8tZ[285], b11_OFWNT9L_8tZ[284], 
        b11_OFWNT9L_8tZ[283], b11_OFWNT9L_8tZ[282], 
        b11_OFWNT9L_8tZ[281], b11_OFWNT9L_8tZ[280], 
        b11_OFWNT9L_8tZ[279], b11_OFWNT9L_8tZ[278], 
        b11_OFWNT9L_8tZ[277], b11_OFWNT9L_8tZ[276], 
        b11_OFWNT9L_8tZ[275], b11_OFWNT9L_8tZ[274], 
        b11_OFWNT9L_8tZ[273], b11_OFWNT9L_8tZ[272], 
        b11_OFWNT9L_8tZ[271], b11_OFWNT9L_8tZ[270], 
        b11_OFWNT9L_8tZ[269], b11_OFWNT9L_8tZ[268], 
        b11_OFWNT9L_8tZ[267], b11_OFWNT9L_8tZ[266], 
        b11_OFWNT9L_8tZ[265], b11_OFWNT9L_8tZ[264], 
        b11_OFWNT9L_8tZ[263], b11_OFWNT9L_8tZ[262], 
        b11_OFWNT9L_8tZ[261], b11_OFWNT9L_8tZ[260], 
        b11_OFWNT9L_8tZ[259], b11_OFWNT9L_8tZ[258], 
        b11_OFWNT9L_8tZ[257], b11_OFWNT9L_8tZ[256], 
        b11_OFWNT9L_8tZ[255], b11_OFWNT9L_8tZ[254], 
        b11_OFWNT9L_8tZ[253], b11_OFWNT9L_8tZ[252], 
        b11_OFWNT9L_8tZ[251], b11_OFWNT9L_8tZ[250], 
        b11_OFWNT9L_8tZ[249], b11_OFWNT9L_8tZ[248], 
        b11_OFWNT9L_8tZ[247], b11_OFWNT9L_8tZ[246], 
        b11_OFWNT9L_8tZ[245], b11_OFWNT9L_8tZ[244], 
        b11_OFWNT9L_8tZ[243], b11_OFWNT9L_8tZ[242], 
        b11_OFWNT9L_8tZ[241], b11_OFWNT9L_8tZ[240], 
        b11_OFWNT9L_8tZ[239], b11_OFWNT9L_8tZ[238], 
        b11_OFWNT9L_8tZ[237], b11_OFWNT9L_8tZ[236], 
        b11_OFWNT9L_8tZ[235], b11_OFWNT9L_8tZ[234], 
        b11_OFWNT9L_8tZ[233], b11_OFWNT9L_8tZ[232], 
        b11_OFWNT9L_8tZ[231], b11_OFWNT9L_8tZ[230], 
        b11_OFWNT9L_8tZ[229], b11_OFWNT9L_8tZ[228], 
        b11_OFWNT9L_8tZ[227], b11_OFWNT9L_8tZ[226], 
        b11_OFWNT9L_8tZ[225], b11_OFWNT9L_8tZ[224], 
        b11_OFWNT9L_8tZ[223], b11_OFWNT9L_8tZ[222], 
        b11_OFWNT9L_8tZ[221], b11_OFWNT9L_8tZ[220], 
        b11_OFWNT9L_8tZ[219], b11_OFWNT9L_8tZ[218], 
        b11_OFWNT9L_8tZ[217], b11_OFWNT9L_8tZ[216], 
        b11_OFWNT9L_8tZ[215], b11_OFWNT9L_8tZ[214], 
        b11_OFWNT9L_8tZ[213], b11_OFWNT9L_8tZ[212], 
        b11_OFWNT9L_8tZ[211], b11_OFWNT9L_8tZ[210], 
        b11_OFWNT9L_8tZ[209], b11_OFWNT9L_8tZ[208], 
        b11_OFWNT9L_8tZ[207], b11_OFWNT9L_8tZ[206], 
        b11_OFWNT9L_8tZ[205], b11_OFWNT9L_8tZ[204], 
        b11_OFWNT9L_8tZ[203], b11_OFWNT9L_8tZ[202], 
        b11_OFWNT9L_8tZ[201], b11_OFWNT9L_8tZ[200], 
        b11_OFWNT9L_8tZ[199], b11_OFWNT9L_8tZ[198], 
        b11_OFWNT9L_8tZ[197], b11_OFWNT9L_8tZ[196], 
        b11_OFWNT9L_8tZ[195], b11_OFWNT9L_8tZ[194], 
        b11_OFWNT9L_8tZ[193], b11_OFWNT9L_8tZ[192], 
        b11_OFWNT9L_8tZ[191], b11_OFWNT9L_8tZ[190], 
        b11_OFWNT9L_8tZ[189], b11_OFWNT9L_8tZ[188], 
        b11_OFWNT9L_8tZ[187], b11_OFWNT9L_8tZ[186], 
        b11_OFWNT9L_8tZ[185], b11_OFWNT9L_8tZ[184], 
        b11_OFWNT9L_8tZ[183], b11_OFWNT9L_8tZ[182], 
        b11_OFWNT9L_8tZ[181], b11_OFWNT9L_8tZ[180], 
        b11_OFWNT9L_8tZ[179], b11_OFWNT9L_8tZ[178], 
        b11_OFWNT9L_8tZ[177], b11_OFWNT9L_8tZ[176], 
        b11_OFWNT9L_8tZ[175], b11_OFWNT9L_8tZ[174], 
        b11_OFWNT9L_8tZ[173], b11_OFWNT9L_8tZ[172], 
        b11_OFWNT9L_8tZ[171], b11_OFWNT9L_8tZ[170], 
        b11_OFWNT9L_8tZ[169], b11_OFWNT9L_8tZ[168], 
        b11_OFWNT9L_8tZ[167], b11_OFWNT9L_8tZ[166], 
        b11_OFWNT9L_8tZ[165], b11_OFWNT9L_8tZ[164], 
        b11_OFWNT9L_8tZ[163], b11_OFWNT9L_8tZ[162], 
        b11_OFWNT9L_8tZ[161], b11_OFWNT9L_8tZ[160], 
        b11_OFWNT9L_8tZ[159], b11_OFWNT9L_8tZ[158], 
        b11_OFWNT9L_8tZ[157], b11_OFWNT9L_8tZ[156], 
        b11_OFWNT9L_8tZ[155], b11_OFWNT9L_8tZ[154], 
        b11_OFWNT9L_8tZ[153], b11_OFWNT9L_8tZ[152], 
        b11_OFWNT9L_8tZ[151], b11_OFWNT9L_8tZ[150], 
        b11_OFWNT9L_8tZ[149], b11_OFWNT9L_8tZ[148], 
        b11_OFWNT9L_8tZ[147], b11_OFWNT9L_8tZ[146], 
        b11_OFWNT9L_8tZ[145], b11_OFWNT9L_8tZ[144], 
        b11_OFWNT9L_8tZ[143], b11_OFWNT9L_8tZ[142], 
        b11_OFWNT9L_8tZ[141], b11_OFWNT9L_8tZ[140], 
        b11_OFWNT9L_8tZ[139], b11_OFWNT9L_8tZ[138], 
        b11_OFWNT9L_8tZ[137], b11_OFWNT9L_8tZ[136], 
        b11_OFWNT9L_8tZ[135], b11_OFWNT9L_8tZ[134], 
        b11_OFWNT9L_8tZ[133], b11_OFWNT9L_8tZ[132], 
        b11_OFWNT9L_8tZ[131], b11_OFWNT9L_8tZ[130], 
        b11_OFWNT9L_8tZ[129], b11_OFWNT9L_8tZ[128], 
        b11_OFWNT9L_8tZ[127], b11_OFWNT9L_8tZ[126], 
        b11_OFWNT9L_8tZ[125], b11_OFWNT9L_8tZ[124], 
        b11_OFWNT9L_8tZ[123], b11_OFWNT9L_8tZ[122], 
        b11_OFWNT9L_8tZ[121], b11_OFWNT9L_8tZ[120], 
        b11_OFWNT9L_8tZ[119], b11_OFWNT9L_8tZ[118], 
        b11_OFWNT9L_8tZ[117], b11_OFWNT9L_8tZ[116], 
        b11_OFWNT9L_8tZ[115], b11_OFWNT9L_8tZ[114], 
        b11_OFWNT9L_8tZ[113], b11_OFWNT9L_8tZ[112], 
        b11_OFWNT9L_8tZ[111], b11_OFWNT9L_8tZ[110], 
        b11_OFWNT9L_8tZ[109], b11_OFWNT9L_8tZ[108], 
        b11_OFWNT9L_8tZ[107], b11_OFWNT9L_8tZ[106], 
        b11_OFWNT9L_8tZ[105], b11_OFWNT9L_8tZ[104], 
        b11_OFWNT9L_8tZ[103], b11_OFWNT9L_8tZ[102], 
        b11_OFWNT9L_8tZ[101], b11_OFWNT9L_8tZ[100], 
        b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], b11_OFWNT9L_8tZ[97], 
        b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], b11_OFWNT9L_8tZ[94], 
        b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], b11_OFWNT9L_8tZ[91], 
        b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], b11_OFWNT9L_8tZ[88], 
        b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], b11_OFWNT9L_8tZ[85], 
        b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], b11_OFWNT9L_8tZ[82], 
        b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], b11_OFWNT9L_8tZ[79], 
        b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], b11_OFWNT9L_8tZ[76], 
        b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], b11_OFWNT9L_8tZ[73], 
        b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], b11_OFWNT9L_8tZ[70], 
        b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], b11_OFWNT9L_8tZ[67], 
        b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], b11_OFWNT9L_8tZ[64], 
        b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], b11_OFWNT9L_8tZ[61], 
        b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], b11_OFWNT9L_8tZ[58], 
        b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], b11_OFWNT9L_8tZ[55], 
        b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], b11_OFWNT9L_8tZ[52], 
        b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], b11_OFWNT9L_8tZ[49], 
        b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], b11_OFWNT9L_8tZ[46], 
        b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], b11_OFWNT9L_8tZ[43], 
        b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], b11_OFWNT9L_8tZ[40], 
        b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], b11_OFWNT9L_8tZ[37], 
        b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], b11_OFWNT9L_8tZ[34], 
        b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], b11_OFWNT9L_8tZ[31], 
        b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], b11_OFWNT9L_8tZ[28], 
        b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], b11_OFWNT9L_8tZ[25], 
        b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], b11_OFWNT9L_8tZ[22], 
        b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], b11_OFWNT9L_8tZ[19], 
        b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], b11_OFWNT9L_8tZ[16], 
        b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], b11_OFWNT9L_8tZ[13], 
        b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], b11_OFWNT9L_8tZ[10], 
        b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], b11_OFWNT9L_8tZ[7], 
        b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], b11_OFWNT9L_8tZ[4], 
        b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], b11_OFWNT9L_8tZ[1], 
        b11_OFWNT9L_8tZ[0]}), .b4_nUAi({\b4_nUAi[1129] , 
        \b4_nUAi[1128] , \b4_nUAi[1127] , \b4_nUAi[1126] , 
        \b4_nUAi[1125] , \b4_nUAi[1124] , \b4_nUAi[1123] , 
        \b4_nUAi[1122] , \b4_nUAi[1121] , \b4_nUAi[1120] , 
        \b4_nUAi[1119] , \b4_nUAi[1118] , \b4_nUAi[1117] , 
        \b4_nUAi[1116] , \b4_nUAi[1115] , \b4_nUAi[1114] , 
        \b4_nUAi[1113] , \b4_nUAi[1112] , \b4_nUAi[1111] , 
        \b4_nUAi[1110] , \b4_nUAi[1109] , \b4_nUAi[1108] , 
        \b4_nUAi[1107] , \b4_nUAi[1106] , \b4_nUAi[1105] , 
        \b4_nUAi[1104] , \b4_nUAi[1103] , \b4_nUAi[1102] , 
        \b4_nUAi[1101] , \b4_nUAi[1100] , \b4_nUAi[1099] , 
        \b4_nUAi[1098] , \b4_nUAi[1097] , \b4_nUAi[1096] , 
        \b4_nUAi[1095] , \b4_nUAi[1094] , \b4_nUAi[1093] , 
        \b4_nUAi[1092] , \b4_nUAi[1091] , \b4_nUAi[1090] , 
        \b4_nUAi[1089] , \b4_nUAi[1088] , \b4_nUAi[1087] , 
        \b4_nUAi[1086] , \b4_nUAi[1085] , \b4_nUAi[1084] , 
        \b4_nUAi[1083] , \b4_nUAi[1082] , \b4_nUAi[1081] , 
        \b4_nUAi[1080] , \b4_nUAi[1079] , \b4_nUAi[1078] , 
        \b4_nUAi[1077] , \b4_nUAi[1076] , \b4_nUAi[1075] , 
        \b4_nUAi[1074] , \b4_nUAi[1073] , \b4_nUAi[1072] , 
        \b4_nUAi[1071] , \b4_nUAi[1070] , \b4_nUAi[1069] , 
        \b4_nUAi[1068] , \b4_nUAi[1067] , \b4_nUAi[1066] , 
        \b4_nUAi[1065] , \b4_nUAi[1064] , \b4_nUAi[1063] , 
        \b4_nUAi[1062] , \b4_nUAi[1061] , \b4_nUAi[1060] , 
        \b4_nUAi[1059] , \b4_nUAi[1058] , \b4_nUAi[1057] , 
        \b4_nUAi[1056] , \b4_nUAi[1055] , \b4_nUAi[1054] , 
        \b4_nUAi[1053] , \b4_nUAi[1052] , \b4_nUAi[1051] , 
        \b4_nUAi[1050] , \b4_nUAi[1049] , \b4_nUAi[1048] , 
        \b4_nUAi[1047] , \b4_nUAi[1046] , \b4_nUAi[1045] , 
        \b4_nUAi[1044] , \b4_nUAi[1043] , \b4_nUAi[1042] , 
        \b4_nUAi[1041] , \b4_nUAi[1040] , \b4_nUAi[1039] , 
        \b4_nUAi[1038] , \b4_nUAi[1037] , \b4_nUAi[1036] , 
        \b4_nUAi[1035] , \b4_nUAi[1034] , \b4_nUAi[1033] , 
        \b4_nUAi[1032] , \b4_nUAi[1031] , \b4_nUAi[1030] , 
        \b4_nUAi[1029] , \b4_nUAi[1028] , \b4_nUAi[1027] , 
        \b4_nUAi[1026] , \b4_nUAi[1025] , \b4_nUAi[1024] , 
        \b4_nUAi[1023] , \b4_nUAi[1022] , \b4_nUAi[1021] , 
        \b4_nUAi[1020] , \b4_nUAi[1019] , \b4_nUAi[1018] , 
        \b4_nUAi[1017] , \b4_nUAi[1016] , \b4_nUAi[1015] , 
        \b4_nUAi[1014] , \b4_nUAi[1013] , \b4_nUAi[1012] , 
        \b4_nUAi[1011] , \b4_nUAi[1010] , \b4_nUAi[1009] , 
        \b4_nUAi[1008] , \b4_nUAi[1007] , \b4_nUAi[1006] , 
        \b4_nUAi[1005] , \b4_nUAi[1004] , \b4_nUAi[1003] , 
        \b4_nUAi[1002] , \b4_nUAi[1001] , \b4_nUAi[1000] , 
        \b4_nUAi[999] , \b4_nUAi[998] , \b4_nUAi[997] , \b4_nUAi[996] , 
        \b4_nUAi[995] , \b4_nUAi[994] , \b4_nUAi[993] , \b4_nUAi[992] , 
        \b4_nUAi[991] , \b4_nUAi[990] , \b4_nUAi[989] , \b4_nUAi[988] , 
        \b4_nUAi[987] , \b4_nUAi[986] , \b4_nUAi[985] , \b4_nUAi[984] , 
        \b4_nUAi[983] , \b4_nUAi[982] , \b4_nUAi[981] , \b4_nUAi[980] , 
        \b4_nUAi[979] , \b4_nUAi[978] , \b4_nUAi[977] , \b4_nUAi[976] , 
        \b4_nUAi[975] , \b4_nUAi[974] , \b4_nUAi[973] , \b4_nUAi[972] , 
        \b4_nUAi[971] , \b4_nUAi[970] , \b4_nUAi[969] , \b4_nUAi[968] , 
        \b4_nUAi[967] , \b4_nUAi[966] , \b4_nUAi[965] , \b4_nUAi[964] , 
        \b4_nUAi[963] , \b4_nUAi[962] , \b4_nUAi[961] , \b4_nUAi[960] , 
        \b4_nUAi[959] , \b4_nUAi[958] , \b4_nUAi[957] , \b4_nUAi[956] , 
        \b4_nUAi[955] , \b4_nUAi[954] , \b4_nUAi[953] , \b4_nUAi[952] , 
        \b4_nUAi[951] , \b4_nUAi[950] , \b4_nUAi[949] , \b4_nUAi[948] , 
        \b4_nUAi[947] , \b4_nUAi[946] , \b4_nUAi[945] , \b4_nUAi[944] , 
        \b4_nUAi[943] , \b4_nUAi[942] , \b4_nUAi[941] , \b4_nUAi[940] , 
        \b4_nUAi[939] , \b4_nUAi[938] , \b4_nUAi[937] , \b4_nUAi[936] , 
        \b4_nUAi[935] , \b4_nUAi[934] , \b4_nUAi[933] , \b4_nUAi[932] , 
        \b4_nUAi[931] , \b4_nUAi[930] , \b4_nUAi[929] , \b4_nUAi[928] , 
        \b4_nUAi[927] , \b4_nUAi[926] , \b4_nUAi[925] , \b4_nUAi[924] , 
        \b4_nUAi[923] , \b4_nUAi[922] , \b4_nUAi[921] , \b4_nUAi[920] , 
        \b4_nUAi[919] , \b4_nUAi[918] , \b4_nUAi[917] , \b4_nUAi[916] , 
        \b4_nUAi[915] , \b4_nUAi[914] , \b4_nUAi[913] , \b4_nUAi[912] , 
        \b4_nUAi[911] , \b4_nUAi[910] , \b4_nUAi[909] , \b4_nUAi[908] , 
        \b4_nUAi[907] , \b4_nUAi[906] , \b4_nUAi[905] , \b4_nUAi[904] , 
        \b4_nUAi[903] , \b4_nUAi[902] , \b4_nUAi[901] , \b4_nUAi[900] , 
        \b4_nUAi[899] , \b4_nUAi[898] , \b4_nUAi[897] , \b4_nUAi[896] , 
        \b4_nUAi[895] , \b4_nUAi[894] , \b4_nUAi[893] , \b4_nUAi[892] , 
        \b4_nUAi[891] , \b4_nUAi[890] , \b4_nUAi[889] , \b4_nUAi[888] , 
        \b4_nUAi[887] , \b4_nUAi[886] , \b4_nUAi[885] , \b4_nUAi[884] , 
        \b4_nUAi[883] , \b4_nUAi[882] , \b4_nUAi[881] , \b4_nUAi[880] , 
        \b4_nUAi[879] , \b4_nUAi[878] , \b4_nUAi[877] , \b4_nUAi[876] , 
        \b4_nUAi[875] , \b4_nUAi[874] , \b4_nUAi[873] , \b4_nUAi[872] , 
        \b4_nUAi[871] , \b4_nUAi[870] , \b4_nUAi[869] , \b4_nUAi[868] , 
        \b4_nUAi[867] , \b4_nUAi[866] , \b4_nUAi[865] , \b4_nUAi[864] , 
        \b4_nUAi[863] , \b4_nUAi[862] , \b4_nUAi[861] , \b4_nUAi[860] , 
        \b4_nUAi[859] , \b4_nUAi[858] , \b4_nUAi[857] , \b4_nUAi[856] , 
        \b4_nUAi[855] , \b4_nUAi[854] , \b4_nUAi[853] , \b4_nUAi[852] , 
        \b4_nUAi[851] , \b4_nUAi[850] , \b4_nUAi[849] , \b4_nUAi[848] , 
        \b4_nUAi[847] , \b4_nUAi[846] , \b4_nUAi[845] , \b4_nUAi[844] , 
        \b4_nUAi[843] , \b4_nUAi[842] , \b4_nUAi[841] , \b4_nUAi[840] , 
        \b4_nUAi[839] , \b4_nUAi[838] , \b4_nUAi[837] , \b4_nUAi[836] , 
        \b4_nUAi[835] , \b4_nUAi[834] , \b4_nUAi[833] , \b4_nUAi[832] , 
        \b4_nUAi[831] , \b4_nUAi[830] , \b4_nUAi[829] , \b4_nUAi[828] , 
        \b4_nUAi[827] , \b4_nUAi[826] , \b4_nUAi[825] , \b4_nUAi[824] , 
        \b4_nUAi[823] , \b4_nUAi[822] , \b4_nUAi[821] , \b4_nUAi[820] , 
        \b4_nUAi[819] , \b4_nUAi[818] , \b4_nUAi[817] , \b4_nUAi[816] , 
        \b4_nUAi[815] , \b4_nUAi[814] , \b4_nUAi[813] , \b4_nUAi[812] , 
        \b4_nUAi[811] , \b4_nUAi[810] , \b4_nUAi[809] , \b4_nUAi[808] , 
        \b4_nUAi[807] , \b4_nUAi[806] , \b4_nUAi[805] , \b4_nUAi[804] , 
        \b4_nUAi[803] , \b4_nUAi[802] , \b4_nUAi[801] , \b4_nUAi[800] , 
        \b4_nUAi[799] , \b4_nUAi[798] , \b4_nUAi[797] , \b4_nUAi[796] , 
        \b4_nUAi[795] , \b4_nUAi[794] , \b4_nUAi[793] , \b4_nUAi[792] , 
        \b4_nUAi[791] , \b4_nUAi[790] , \b4_nUAi[789] , \b4_nUAi[788] , 
        \b4_nUAi[787] , \b4_nUAi[786] , \b4_nUAi[785] , \b4_nUAi[784] , 
        \b4_nUAi[783] , \b4_nUAi[782] , \b4_nUAi[781] , \b4_nUAi[780] , 
        \b4_nUAi[779] , \b4_nUAi[778] , \b4_nUAi[777] , \b4_nUAi[776] , 
        \b4_nUAi[775] , \b4_nUAi[774] , \b4_nUAi[773] , \b4_nUAi[772] , 
        \b4_nUAi[771] , \b4_nUAi[770] , \b4_nUAi[769] , \b4_nUAi[768] , 
        \b4_nUAi[767] , \b4_nUAi[766] , \b4_nUAi[765] , \b4_nUAi[764] , 
        \b4_nUAi[763] , \b4_nUAi[762] , \b4_nUAi[761] , \b4_nUAi[760] , 
        \b4_nUAi[759] , \b4_nUAi[758] , \b4_nUAi[757] , \b4_nUAi[756] , 
        \b4_nUAi[755] , \b4_nUAi[754] , \b4_nUAi[753] , \b4_nUAi[752] , 
        \b4_nUAi[751] , \b4_nUAi[750] , \b4_nUAi[749] , \b4_nUAi[748] , 
        \b4_nUAi[747] , \b4_nUAi[746] , \b4_nUAi[745] , \b4_nUAi[744] , 
        \b4_nUAi[743] , \b4_nUAi[742] , \b4_nUAi[741] , \b4_nUAi[740] , 
        \b4_nUAi[739] , \b4_nUAi[738] , \b4_nUAi[737] , \b4_nUAi[736] , 
        \b4_nUAi[735] , \b4_nUAi[734] , \b4_nUAi[733] , \b4_nUAi[732] , 
        \b4_nUAi[731] , \b4_nUAi[730] , \b4_nUAi[729] , \b4_nUAi[728] , 
        \b4_nUAi[727] , \b4_nUAi[726] , \b4_nUAi[725] , \b4_nUAi[724] , 
        \b4_nUAi[723] , \b4_nUAi[722] , \b4_nUAi[721] , \b4_nUAi[720] , 
        \b4_nUAi[719] , \b4_nUAi[718] , \b4_nUAi[717] , \b4_nUAi[716] , 
        \b4_nUAi[715] , \b4_nUAi[714] , \b4_nUAi[713] , \b4_nUAi[712] , 
        \b4_nUAi[711] , \b4_nUAi[710] , \b4_nUAi[709] , \b4_nUAi[708] , 
        \b4_nUAi[707] , \b4_nUAi[706] , \b4_nUAi[705] , \b4_nUAi[704] , 
        \b4_nUAi[703] , \b4_nUAi[702] , \b4_nUAi[701] , \b4_nUAi[700] , 
        \b4_nUAi[699] , \b4_nUAi[698] , \b4_nUAi[697] , \b4_nUAi[696] , 
        \b4_nUAi[695] , \b4_nUAi[694] , \b4_nUAi[693] , \b4_nUAi[692] , 
        \b4_nUAi[691] , \b4_nUAi[690] , \b4_nUAi[689] , \b4_nUAi[688] , 
        \b4_nUAi[687] , \b4_nUAi[686] , \b4_nUAi[685] , \b4_nUAi[684] , 
        \b4_nUAi[683] , \b4_nUAi[682] , \b4_nUAi[681] , \b4_nUAi[680] , 
        \b4_nUAi[679] , \b4_nUAi[678] , \b4_nUAi[677] , \b4_nUAi[676] , 
        \b4_nUAi[675] , \b4_nUAi[674] , \b4_nUAi[673] , \b4_nUAi[672] , 
        \b4_nUAi[671] , \b4_nUAi[670] , \b4_nUAi[669] , \b4_nUAi[668] , 
        \b4_nUAi[667] , \b4_nUAi[666] , \b4_nUAi[665] , \b4_nUAi[664] , 
        \b4_nUAi[663] , \b4_nUAi[662] , \b4_nUAi[661] , \b4_nUAi[660] , 
        \b4_nUAi[659] , \b4_nUAi[658] , \b4_nUAi[657] , \b4_nUAi[656] , 
        \b4_nUAi[655] , \b4_nUAi[654] , \b4_nUAi[653] , \b4_nUAi[652] , 
        \b4_nUAi[651] , \b4_nUAi[650] , \b4_nUAi[649] , \b4_nUAi[648] , 
        \b4_nUAi[647] , \b4_nUAi[646] , \b4_nUAi[645] , \b4_nUAi[644] , 
        \b4_nUAi[643] , \b4_nUAi[642] , \b4_nUAi[641] , \b4_nUAi[640] , 
        \b4_nUAi[639] , \b4_nUAi[638] , \b4_nUAi[637] , \b4_nUAi[636] , 
        \b4_nUAi[635] , \b4_nUAi[634] , \b4_nUAi[633] , \b4_nUAi[632] , 
        \b4_nUAi[631] , \b4_nUAi[630] , \b4_nUAi[629] , \b4_nUAi[628] , 
        \b4_nUAi[627] , \b4_nUAi[626] , \b4_nUAi[625] , \b4_nUAi[624] , 
        \b4_nUAi[623] , \b4_nUAi[622] , \b4_nUAi[621] , \b4_nUAi[620] , 
        \b4_nUAi[619] , \b4_nUAi[618] , \b4_nUAi[617] , \b4_nUAi[616] , 
        \b4_nUAi[615] , \b4_nUAi[614] , \b4_nUAi[613] , \b4_nUAi[612] , 
        \b4_nUAi[611] , \b4_nUAi[610] , \b4_nUAi[609] , \b4_nUAi[608] , 
        \b4_nUAi[607] , \b4_nUAi[606] , \b4_nUAi[605] , \b4_nUAi[604] , 
        \b4_nUAi[603] , \b4_nUAi[602] , \b4_nUAi[601] , \b4_nUAi[600] , 
        \b4_nUAi[599] , \b4_nUAi[598] , \b4_nUAi[597] , \b4_nUAi[596] , 
        \b4_nUAi[595] , \b4_nUAi[594] , \b4_nUAi[593] , \b4_nUAi[592] , 
        \b4_nUAi[591] , \b4_nUAi[590] , \b4_nUAi[589] , \b4_nUAi[588] , 
        \b4_nUAi[587] , \b4_nUAi[586] , \b4_nUAi[585] , \b4_nUAi[584] , 
        \b4_nUAi[583] , \b4_nUAi[582] , \b4_nUAi[581] , \b4_nUAi[580] , 
        \b4_nUAi[579] , \b4_nUAi[578] , \b4_nUAi[577] , \b4_nUAi[576] , 
        \b4_nUAi[575] , \b4_nUAi[574] , \b4_nUAi[573] , \b4_nUAi[572] , 
        \b4_nUAi[571] , \b4_nUAi[570] , \b4_nUAi[569] , \b4_nUAi[568] , 
        \b4_nUAi[567] , \b4_nUAi[566] , \b4_nUAi[565] , \b4_nUAi[564] , 
        \b4_nUAi[563] , \b4_nUAi[562] , \b4_nUAi[561] , \b4_nUAi[560] , 
        \b4_nUAi[559] , \b4_nUAi[558] , \b4_nUAi[557] , \b4_nUAi[556] , 
        \b4_nUAi[555] , \b4_nUAi[554] , \b4_nUAi[553] , \b4_nUAi[552] , 
        \b4_nUAi[551] , \b4_nUAi[550] , \b4_nUAi[549] , \b4_nUAi[548] , 
        \b4_nUAi[547] , \b4_nUAi[546] , \b4_nUAi[545] , \b4_nUAi[544] , 
        \b4_nUAi[543] , \b4_nUAi[542] , \b4_nUAi[541] , \b4_nUAi[540] , 
        \b4_nUAi[539] , \b4_nUAi[538] , \b4_nUAi[537] , \b4_nUAi[536] , 
        \b4_nUAi[535] , \b4_nUAi[534] , \b4_nUAi[533] , \b4_nUAi[532] , 
        \b4_nUAi[531] , \b4_nUAi[530] , \b4_nUAi[529] , \b4_nUAi[528] , 
        \b4_nUAi[527] , \b4_nUAi[526] , \b4_nUAi[525] , \b4_nUAi[524] , 
        \b4_nUAi[523] , \b4_nUAi[522] , \b4_nUAi[521] , \b4_nUAi[520] , 
        \b4_nUAi[519] , \b4_nUAi[518] , \b4_nUAi[517] , \b4_nUAi[516] , 
        \b4_nUAi[515] , \b4_nUAi[514] , \b4_nUAi[513] , \b4_nUAi[512] , 
        \b4_nUAi[511] , \b4_nUAi[510] , \b4_nUAi[509] , \b4_nUAi[508] , 
        \b4_nUAi[507] , \b4_nUAi[506] , \b4_nUAi[505] , \b4_nUAi[504] , 
        \b4_nUAi[503] , \b4_nUAi[502] , \b4_nUAi[501] , \b4_nUAi[500] , 
        \b4_nUAi[499] , \b4_nUAi[498] , \b4_nUAi[497] , \b4_nUAi[496] , 
        \b4_nUAi[495] , \b4_nUAi[494] , \b4_nUAi[493] , \b4_nUAi[492] , 
        \b4_nUAi[491] , \b4_nUAi[490] , \b4_nUAi[489] , \b4_nUAi[488] , 
        \b4_nUAi[487] , \b4_nUAi[486] , \b4_nUAi[485] , \b4_nUAi[484] , 
        \b4_nUAi[483] , \b4_nUAi[482] , \b4_nUAi[481] , \b4_nUAi[480] , 
        \b4_nUAi[479] , \b4_nUAi[478] , \b4_nUAi[477] , \b4_nUAi[476] , 
        \b4_nUAi[475] , \b4_nUAi[474] , \b4_nUAi[473] , \b4_nUAi[472] , 
        \b4_nUAi[471] , \b4_nUAi[470] , \b4_nUAi[469] , \b4_nUAi[468] , 
        \b4_nUAi[467] , \b4_nUAi[466] , \b4_nUAi[465] , \b4_nUAi[464] , 
        \b4_nUAi[463] , \b4_nUAi[462] , \b4_nUAi[461] , \b4_nUAi[460] , 
        \b4_nUAi[459] , \b4_nUAi[458] , \b4_nUAi[457] , \b4_nUAi[456] , 
        \b4_nUAi[455] , \b4_nUAi[454] , \b4_nUAi[453] , \b4_nUAi[452] , 
        \b4_nUAi[451] , \b4_nUAi[450] , \b4_nUAi[449] , \b4_nUAi[448] , 
        \b4_nUAi[447] , \b4_nUAi[446] , \b4_nUAi[445] , \b4_nUAi[444] , 
        \b4_nUAi[443] , \b4_nUAi[442] , \b4_nUAi[441] , \b4_nUAi[440] , 
        \b4_nUAi[439] , \b4_nUAi[438] , \b4_nUAi[437] , \b4_nUAi[436] , 
        \b4_nUAi[435] , \b4_nUAi[434] , \b4_nUAi[433] , \b4_nUAi[432] , 
        \b4_nUAi[431] , \b4_nUAi[430] , \b4_nUAi[429] , \b4_nUAi[428] , 
        \b4_nUAi[427] , \b4_nUAi[426] , \b4_nUAi[425] , \b4_nUAi[424] , 
        \b4_nUAi[423] , \b4_nUAi[422] , \b4_nUAi[421] , \b4_nUAi[420] , 
        \b4_nUAi[419] , \b4_nUAi[418] , \b4_nUAi[417] , \b4_nUAi[416] , 
        \b4_nUAi[415] , \b4_nUAi[414] , \b4_nUAi[413] , \b4_nUAi[412] , 
        \b4_nUAi[411] , \b4_nUAi[410] , \b4_nUAi[409] , \b4_nUAi[408] , 
        \b4_nUAi[407] , \b4_nUAi[406] , \b4_nUAi[405] , \b4_nUAi[404] , 
        \b4_nUAi[403] , \b4_nUAi[402] , \b4_nUAi[401] , \b4_nUAi[400] , 
        \b4_nUAi[399] , \b4_nUAi[398] , \b4_nUAi[397] , \b4_nUAi[396] , 
        \b4_nUAi[395] , \b4_nUAi[394] , \b4_nUAi[393] , \b4_nUAi[392] , 
        \b4_nUAi[391] , \b4_nUAi[390] , \b4_nUAi[389] , \b4_nUAi[388] , 
        \b4_nUAi[387] , \b4_nUAi[386] , \b4_nUAi[385] , \b4_nUAi[384] , 
        \b4_nUAi[383] , \b4_nUAi[382] , \b4_nUAi[381] , \b4_nUAi[380] , 
        \b4_nUAi[379] , \b4_nUAi[378] , \b4_nUAi[377] , \b4_nUAi[376] , 
        \b4_nUAi[375] , \b4_nUAi[374] , \b4_nUAi[373] , \b4_nUAi[372] , 
        \b4_nUAi[371] , \b4_nUAi[370] , \b4_nUAi[369] , \b4_nUAi[368] , 
        \b4_nUAi[367] , \b4_nUAi[366] , \b4_nUAi[365] , \b4_nUAi[364] , 
        \b4_nUAi[363] , \b4_nUAi[362] , \b4_nUAi[361] , \b4_nUAi[360] , 
        \b4_nUAi[359] , \b4_nUAi[358] , \b4_nUAi[357] , \b4_nUAi[356] , 
        \b4_nUAi[355] , \b4_nUAi[354] , \b4_nUAi[353] , \b4_nUAi[352] , 
        \b4_nUAi[351] , \b4_nUAi[350] , \b4_nUAi[349] , \b4_nUAi[348] , 
        \b4_nUAi[347] , \b4_nUAi[346] , \b4_nUAi[345] , \b4_nUAi[344] , 
        \b4_nUAi[343] , \b4_nUAi[342] , \b4_nUAi[341] , \b4_nUAi[340] , 
        \b4_nUAi[339] , \b4_nUAi[338] , \b4_nUAi[337] , \b4_nUAi[336] , 
        \b4_nUAi[335] , \b4_nUAi[334] , \b4_nUAi[333] , \b4_nUAi[332] , 
        \b4_nUAi[331] , \b4_nUAi[330] , \b4_nUAi[329] , \b4_nUAi[328] , 
        \b4_nUAi[327] , \b4_nUAi[326] , \b4_nUAi[325] , \b4_nUAi[324] , 
        \b4_nUAi[323] , \b4_nUAi[322] , \b4_nUAi[321] , \b4_nUAi[320] , 
        \b4_nUAi[319] , \b4_nUAi[318] , \b4_nUAi[317] , \b4_nUAi[316] , 
        \b4_nUAi[315] , \b4_nUAi[314] , \b4_nUAi[313] , \b4_nUAi[312] , 
        \b4_nUAi[311] , \b4_nUAi[310] , \b4_nUAi[309] , \b4_nUAi[308] , 
        \b4_nUAi[307] , \b4_nUAi[306] , \b4_nUAi[305] , \b4_nUAi[304] , 
        \b4_nUAi[303] , \b4_nUAi[302] , \b4_nUAi[301] , \b4_nUAi[300] , 
        \b4_nUAi[299] , \b4_nUAi[298] , \b4_nUAi[297] , \b4_nUAi[296] , 
        \b4_nUAi[295] , \b4_nUAi[294] , \b4_nUAi[293] , \b4_nUAi[292] , 
        \b4_nUAi[291] , \b4_nUAi[290] , \b4_nUAi[289] , \b4_nUAi[288] , 
        \b4_nUAi[287] , \b4_nUAi[286] , \b4_nUAi[285] , \b4_nUAi[284] , 
        \b4_nUAi[283] , \b4_nUAi[282] , \b4_nUAi[281] , \b4_nUAi[280] , 
        \b4_nUAi[279] , \b4_nUAi[278] , \b4_nUAi[277] , \b4_nUAi[276] , 
        \b4_nUAi[275] , \b4_nUAi[274] , \b4_nUAi[273] , \b4_nUAi[272] , 
        \b4_nUAi[271] , \b4_nUAi[270] , \b4_nUAi[269] , \b4_nUAi[268] , 
        \b4_nUAi[267] , \b4_nUAi[266] , \b4_nUAi[265] , \b4_nUAi[264] , 
        \b4_nUAi[263] , \b4_nUAi[262] , \b4_nUAi[261] , \b4_nUAi[260] , 
        \b4_nUAi[259] , \b4_nUAi[258] , \b4_nUAi[257] , \b4_nUAi[256] , 
        \b4_nUAi[255] , \b4_nUAi[254] , \b4_nUAi[253] , \b4_nUAi[252] , 
        \b4_nUAi[251] , \b4_nUAi[250] , \b4_nUAi[249] , \b4_nUAi[248] , 
        \b4_nUAi[247] , \b4_nUAi[246] , \b4_nUAi[245] , \b4_nUAi[244] , 
        \b4_nUAi[243] , \b4_nUAi[242] , \b4_nUAi[241] , \b4_nUAi[240] , 
        \b4_nUAi[239] , \b4_nUAi[238] , \b4_nUAi[237] , \b4_nUAi[236] , 
        \b4_nUAi[235] , \b4_nUAi[234] , \b4_nUAi[233] , \b4_nUAi[232] , 
        \b4_nUAi[231] , \b4_nUAi[230] , \b4_nUAi[229] , \b4_nUAi[228] , 
        \b4_nUAi[227] , \b4_nUAi[226] , \b4_nUAi[225] , \b4_nUAi[224] , 
        \b4_nUAi[223] , \b4_nUAi[222] , \b4_nUAi[221] , \b4_nUAi[220] , 
        \b4_nUAi[219] , \b4_nUAi[218] , \b4_nUAi[217] , \b4_nUAi[216] , 
        \b4_nUAi[215] , \b4_nUAi[214] , \b4_nUAi[213] , \b4_nUAi[212] , 
        \b4_nUAi[211] , \b4_nUAi[210] , \b4_nUAi[209] , \b4_nUAi[208] , 
        \b4_nUAi[207] , \b4_nUAi[206] , \b4_nUAi[205] , \b4_nUAi[204] , 
        \b4_nUAi[203] , \b4_nUAi[202] , \b4_nUAi[201] , \b4_nUAi[200] , 
        \b4_nUAi[199] , \b4_nUAi[198] , \b4_nUAi[197] , \b4_nUAi[196] , 
        \b4_nUAi[195] , \b4_nUAi[194] , \b4_nUAi[193] , \b4_nUAi[192] , 
        \b4_nUAi[191] , \b4_nUAi[190] , \b4_nUAi[189] , \b4_nUAi[188] , 
        \b4_nUAi[187] , \b4_nUAi[186] , \b4_nUAi[185] , \b4_nUAi[184] , 
        \b4_nUAi[183] , \b4_nUAi[182] , \b4_nUAi[181] , \b4_nUAi[180] , 
        \b4_nUAi[179] , \b4_nUAi[178] , \b4_nUAi[177] , \b4_nUAi[176] , 
        \b4_nUAi[175] , \b4_nUAi[174] , \b4_nUAi[173] , \b4_nUAi[172] , 
        \b4_nUAi[171] , \b4_nUAi[170] , \b4_nUAi[169] , \b4_nUAi[168] , 
        \b4_nUAi[167] , \b4_nUAi[166] , \b4_nUAi[165] , \b4_nUAi[164] , 
        \b4_nUAi[163] , \b4_nUAi[162] , \b4_nUAi[161] , \b4_nUAi[160] , 
        \b4_nUAi[159] , \b4_nUAi[158] , \b4_nUAi[157] , \b4_nUAi[156] , 
        \b4_nUAi[155] , \b4_nUAi[154] , \b4_nUAi[153] , \b4_nUAi[152] , 
        \b4_nUAi[151] , \b4_nUAi[150] , \b4_nUAi[149] , \b4_nUAi[148] , 
        \b4_nUAi[147] , \b4_nUAi[146] , \b4_nUAi[145] , \b4_nUAi[144] , 
        \b4_nUAi[143] , \b4_nUAi[142] , \b4_nUAi[141] , \b4_nUAi[140] , 
        \b4_nUAi[139] , \b4_nUAi[138] , \b4_nUAi[137] , \b4_nUAi[136] , 
        \b4_nUAi[135] , \b4_nUAi[134] , \b4_nUAi[133] , \b4_nUAi[132] , 
        \b4_nUAi[131] , \b4_nUAi[130] , \b4_nUAi[129] , \b4_nUAi[128] , 
        \b4_nUAi[127] , \b4_nUAi[126] , \b4_nUAi[125] , \b4_nUAi[124] , 
        \b4_nUAi[123] , \b4_nUAi[122] , \b4_nUAi[121] , \b4_nUAi[120] , 
        \b4_nUAi[119] , \b4_nUAi[118] , \b4_nUAi[117] , \b4_nUAi[116] , 
        \b4_nUAi[115] , \b4_nUAi[114] , \b4_nUAi[113] , \b4_nUAi[112] , 
        \b4_nUAi[111] , \b4_nUAi[110] , \b4_nUAi[109] , \b4_nUAi[108] , 
        \b4_nUAi[107] , \b4_nUAi[106] , \b4_nUAi[105] , \b4_nUAi[104] , 
        \b4_nUAi[103] , \b4_nUAi[102] , \b4_nUAi[101] , \b4_nUAi[100] , 
        \b4_nUAi[99] , \b4_nUAi[98] , \b4_nUAi[97] , \b4_nUAi[96] , 
        \b4_nUAi[95] , \b4_nUAi[94] , \b4_nUAi[93] , \b4_nUAi[92] , 
        \b4_nUAi[91] , \b4_nUAi[90] , \b4_nUAi[89] , \b4_nUAi[88] , 
        \b4_nUAi[87] , \b4_nUAi[86] , \b4_nUAi[85] , \b4_nUAi[84] , 
        \b4_nUAi[83] , \b4_nUAi[82] , \b4_nUAi[81] , \b4_nUAi[80] , 
        \b4_nUAi[79] , \b4_nUAi[78] , \b4_nUAi[77] , \b4_nUAi[76] , 
        \b4_nUAi[75] , \b4_nUAi[74] , \b4_nUAi[73] , \b4_nUAi[72] , 
        \b4_nUAi[71] , \b4_nUAi[70] , \b4_nUAi[69] , \b4_nUAi[68] , 
        \b4_nUAi[67] , \b4_nUAi[66] , \b4_nUAi[65] , \b4_nUAi[64] , 
        \b4_nUAi[63] , \b4_nUAi[62] , \b4_nUAi[61] , \b4_nUAi[60] , 
        \b4_nUAi[59] , \b4_nUAi[58] , \b4_nUAi[57] , \b4_nUAi[56] , 
        \b4_nUAi[55] , \b4_nUAi[54] , \b4_nUAi[53] , \b4_nUAi[52] , 
        \b4_nUAi[51] , \b4_nUAi[50] , \b4_nUAi[49] , \b4_nUAi[48] , 
        \b4_nUAi[47] , \b4_nUAi[46] , \b4_nUAi[45] , \b4_nUAi[44] , 
        \b4_nUAi[43] , \b4_nUAi[42] , \b4_nUAi[41] , \b4_nUAi[40] , 
        \b4_nUAi[39] , \b4_nUAi[38] , \b4_nUAi[37] , \b4_nUAi[36] , 
        \b4_nUAi[35] , \b4_nUAi[34] , \b4_nUAi[33] , \b4_nUAi[32] , 
        \b4_nUAi[31] , \b4_nUAi[30] , \b4_nUAi[29] , \b4_nUAi[28] , 
        \b4_nUAi[27] , \b4_nUAi[26] , \b4_nUAi[25] , \b4_nUAi[24] , 
        \b4_nUAi[23] , \b4_nUAi[22] , \b4_nUAi[21] , \b4_nUAi[20] , 
        \b4_nUAi[19] , \b4_nUAi[18] , \b4_nUAi[17] , \b4_nUAi[16] , 
        \b4_nUAi[15] , \b4_nUAi[14] , \b4_nUAi[13] , \b4_nUAi[12] , 
        \b4_nUAi[11] , \b4_nUAi[10] , \b4_nUAi[9] , \b4_nUAi[8] , 
        \b4_nUAi[7] , \b4_nUAi[6] , \b4_nUAi[5] , \b4_nUAi[4] , 
        \b4_nUAi[3] , \b4_nUAi[2] , \b4_nUAi[1] , \b4_nUAi[0] }), 
        .b11_uUT0JC4gFrY({\b11_uUT0JC4gFrY[1] }), .BW_clk_c(BW_clk_c), 
        .b7_PSyi3wy(b7_PSyi3wy));
    GND GND (.Y(GND_net_1));
    SLE b7_PSyil9s (.D(\b11_uUT0JC4gFrY[1] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b11_PSyil9s_FMZ));
    
endmodule


module b8_nR_ymqrG_10s_5s_0_0s_0s_1_510_x_0(
       b6_nfs_IF_i_0,
       b6_nUT_IF,
       b6_nfs_IF,
       IICE_comm2iice_3,
       IICE_comm2iice_0,
       IICE_comm2iice_2,
       b4_PLyF,
       b13_nUTQBgfDb_Z4D,
       b12_nUTQBgfDb_bd,
       b16_nYhI39swMeEd_A78,
       b15_nYhI39swMeEd_Mg,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_qH,
       b11_vABZ3qsY_XH
    );
output [1:1] b6_nfs_IF_i_0;
output [9:0] b6_nUT_IF;
output [4:0] b6_nfs_IF;
input  IICE_comm2iice_3;
input  IICE_comm2iice_0;
input  IICE_comm2iice_2;
input  b4_PLyF;
output b13_nUTQBgfDb_Z4D;
input  b12_nUTQBgfDb_bd;
output b16_nYhI39swMeEd_A78;
input  b15_nYhI39swMeEd_Mg;
output b12_vABZ3qsY_Lyh;
output b11_vABZ3qsY_qH;
input  b11_vABZ3qsY_XH;

    wire \b10_nUT_M9kYfr[2]_net_1 , VCC_net_1, 
        \b10_nUT_M9kYfr[3]_net_1 , b10_nUT_M9kYfr4_net_1, GND_net_1, 
        \b10_nUT_M9kYfr[4]_net_1 , \b10_nUT_M9kYfr[5]_net_1 , 
        \b10_nUT_M9kYfr[6]_net_1 , \b10_nUT_M9kYfr[7]_net_1 , 
        \b10_nUT_M9kYfr[8]_net_1 , \b10_nUT_M9kYfr[9]_net_1 , 
        \b10_nfs_M9kYfr[1]_net_1 , b10_nfs_M9kYfr4_net_1, 
        \b10_nfs_M9kYfr[2]_net_1 , \b10_nfs_M9kYfr[3]_net_1 , 
        \b10_nfs_M9kYfr[4]_net_1 , \b10_nUT_M9kYfr[1]_net_1 , 
        b15_vABZ3qsY_ub3Rme3_net_1, b8_vABZ3qsY_RNO;
    
    SLE \genblk1.b3_nfs[4]  (.D(\b10_nfs_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[4]));
    SLE \b10_nUT_M9kYfr[6]  (.D(\b10_nUT_M9kYfr[7]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[6]_net_1 ));
    SLE \genblk2.b3_nUT[9]  (.D(\b10_nUT_M9kYfr[9]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[9]));
    CFG1 #( .INIT(2'h1) )  \genblk1.b3_nfs_RNI8HD5[1]  (.A(
        b6_nfs_IF[1]), .Y(b6_nfs_IF_i_0[1]));
    SLE \genblk2.b3_nUT[6]  (.D(\b10_nUT_M9kYfr[6]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[6]));
    SLE \b10_nUT_M9kYfr[9]  (.D(b4_PLyF), .CLK(IICE_comm2iice_3), .EN(
        b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b10_nUT_M9kYfr[9]_net_1 ));
    CFG2 #( .INIT(4'h8) )  b10_nfs_M9kYfr4 (.A(b12_nUTQBgfDb_bd), .B(
        IICE_comm2iice_2), .Y(b10_nfs_M9kYfr4_net_1));
    SLE \genblk2.b3_nUT[3]  (.D(\b10_nUT_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[3]));
    SLE \b10_nfs_M9kYfr[2]  (.D(\b10_nfs_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nfs_M9kYfr[2]_net_1 ));
    SLE \genblk2.b3_nUT[2]  (.D(\b10_nUT_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[2]));
    SLE \b10_nUT_M9kYfr[3]  (.D(\b10_nUT_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[3]_net_1 ));
    SLE b15_vABZ3qsY_ub3Rme (.D(b4_PLyF), .CLK(IICE_comm2iice_3), .EN(
        b15_vABZ3qsY_ub3Rme3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b12_vABZ3qsY_Lyh));
    VCC VCC (.Y(VCC_net_1));
    SLE \b10_nfs_M9kYfr[3]  (.D(\b10_nfs_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nfs_M9kYfr[3]_net_1 ));
    SLE \genblk1.b3_nfs[3]  (.D(\b10_nfs_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[3]));
    SLE \genblk2.b3_nUT[7]  (.D(\b10_nUT_M9kYfr[7]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[7]));
    SLE \genblk1.b3_nfs[1]  (.D(\b10_nfs_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[1]));
    SLE \b10_nfs_M9kYfr[1]  (.D(\b10_nfs_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nfs_M9kYfr[1]_net_1 ));
    SLE \b10_nUT_M9kYfr[4]  (.D(\b10_nUT_M9kYfr[5]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[4]_net_1 ));
    SLE \genblk2.b3_nUT[0]  (.D(b16_nYhI39swMeEd_A78), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[0]));
    SLE \b10_nUT_M9kYfr[1]  (.D(\b10_nUT_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[1]_net_1 ));
    SLE \b10_nUT_M9kYfr[0]  (.D(\b10_nUT_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b16_nYhI39swMeEd_A78));
    GND GND (.Y(GND_net_1));
    SLE \genblk2.b3_nUT[8]  (.D(\b10_nUT_M9kYfr[8]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[8]));
    SLE \b10_nfs_M9kYfr[4]  (.D(b4_PLyF), .CLK(IICE_comm2iice_3), .EN(
        b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b10_nfs_M9kYfr[4]_net_1 ));
    SLE \genblk2.b3_nUT[4]  (.D(\b10_nUT_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[4]));
    SLE \b10_nfs_M9kYfr[0]  (.D(\b10_nfs_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b13_nUTQBgfDb_Z4D));
    SLE \b10_nUT_M9kYfr[7]  (.D(\b10_nUT_M9kYfr[8]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  b10_nUT_M9kYfr4 (.A(b15_nYhI39swMeEd_Mg), 
        .B(IICE_comm2iice_2), .Y(b10_nUT_M9kYfr4_net_1));
    SLE \b10_nUT_M9kYfr[8]  (.D(\b10_nUT_M9kYfr[9]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[8]_net_1 ));
    SLE \genblk1.b3_nfs[2]  (.D(\b10_nfs_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[2]));
    SLE \genblk1.b3_nfs[0]  (.D(b13_nUTQBgfDb_Z4D), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[0]));
    SLE \genblk3.b8_vABZ3qsY  (.D(b12_vABZ3qsY_Lyh), .CLK(
        IICE_comm2iice_0), .EN(b8_vABZ3qsY_RNO), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b11_vABZ3qsY_qH));
    SLE \b10_nUT_M9kYfr[5]  (.D(\b10_nUT_M9kYfr[6]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[5]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \genblk3.b8_vABZ3qsY_RNO  (.A(
        b11_vABZ3qsY_XH), .B(b6_nfs_IF[1]), .Y(b8_vABZ3qsY_RNO));
    SLE \genblk2.b3_nUT[5]  (.D(\b10_nUT_M9kYfr[5]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[5]));
    CFG2 #( .INIT(4'h8) )  b15_vABZ3qsY_ub3Rme3 (.A(b11_vABZ3qsY_XH), 
        .B(IICE_comm2iice_2), .Y(b15_vABZ3qsY_ub3Rme3_net_1));
    SLE \b10_nUT_M9kYfr[2]  (.D(\b10_nUT_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[2]_net_1 ));
    SLE \genblk2.b3_nUT[1]  (.D(\b10_nUT_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[1]));
    
endmodule


module clock2_en_reg_en_5s_x_0(
       IICE_comm2iice,
       b6_nfs_IF_i_0,
       status_b2sclk,
       b6_nfs_IF,
       b6_Ocm0rW,
       b6_Ocm0rW_0_i_a2_1,
       b13_nAzGfFM_sLsv3_3,
       b13_nAzGfFM_sLsv3_0,
       b13_nAzGfFM_sLsv3_2,
       BW_clk_c,
       N_38
    );
input  [11:11] IICE_comm2iice;
input  [1:1] b6_nfs_IF_i_0;
output [3:0] status_b2sclk;
input  [1:1] b6_nfs_IF;
input  [2:2] b6_Ocm0rW;
input  [1:1] b6_Ocm0rW_0_i_a2_1;
input  b13_nAzGfFM_sLsv3_3;
input  b13_nAzGfFM_sLsv3_0;
input  b13_nAzGfFM_sLsv3_2;
input  BW_clk_c;
input  N_38;

    wire src_ack_net_1, src_ack_i_0, VCC_net_1, \int_data[0]_net_1 , 
        dout4_0_a2_RNIKLH5_net_1, GND_net_1, \int_data[1]_net_1 , 
        \int_data[2]_net_1 , \int_data[3]_net_1 , dout4, N_148_i_0, 
        in_en_RNICUKI_net_1, N_19_i_0, in_en_net_1, src_req_net_1, 
        src_req_RNO_0_net_1, in_enc_1_i, N_156_i_0, in_enc_net_1, 
        dst_req_d_net_1, dst_req_d_0, dst_req_net_1, dst_req_0;
    
    SLE \dout[1]  (.D(\int_data[1]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[1]));
    CFG2 #( .INIT(4'h4) )  dst_req_r (.A(b6_nfs_IF[1]), .B(
        src_req_net_1), .Y(dst_req_0));
    CFG2 #( .INIT(4'hE) )  src_req_RNO_0 (.A(in_enc_1_i), .B(
        b6_nfs_IF[1]), .Y(src_req_RNO_0_net_1));
    CFG3 #( .INIT(8'hAB) )  \int_data_RNO[1]  (.A(b13_nAzGfFM_sLsv3_2), 
        .B(b6_Ocm0rW_0_i_a2_1[1]), .C(N_38), .Y(N_19_i_0));
    SLE \dout[3]  (.D(\int_data[3]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[3]));
    SLE \int_data[1]  (.D(N_19_i_0), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[1]_net_1 ));
    SLE \dout[2]  (.D(\int_data[2]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[2]));
    GND GND (.Y(GND_net_1));
    SLE in_en (.D(in_enc_net_1), .CLK(BW_clk_c), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(b6_nfs_IF_i_0[1]), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(in_en_net_1));
    CFG2 #( .INIT(4'hE) )  src_ack_RNO (.A(dst_req_net_1), .B(
        dst_req_d_net_1), .Y(N_156_i_0));
    SLE src_ack (.D(N_156_i_0), .CLK(BW_clk_c), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(b6_nfs_IF_i_0[1]), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(src_ack_net_1));
    SLE \int_data[0]  (.D(N_148_i_0), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[0]_net_1 ));
    SLE \int_data[2]  (.D(b6_Ocm0rW[2]), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[2]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \int_data_RNO[0]  (.A(N_38), .B(
        b13_nAzGfFM_sLsv3_0), .Y(N_148_i_0));
    SLE \dout[0]  (.D(\int_data[0]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[0]));
    CFG2 #( .INIT(4'hE) )  src_req_RNO_1 (.A(in_en_net_1), .B(
        src_ack_net_1), .Y(in_enc_1_i));
    CFG3 #( .INIT(8'h01) )  in_enc (.A(src_req_net_1), .B(
        src_ack_net_1), .C(in_en_net_1), .Y(in_enc_net_1));
    SLE dst_req (.D(dst_req_0), .CLK(IICE_comm2iice[11]), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dst_req_net_1));
    CFG1 #( .INIT(2'h1) )  src_req_RNO (.A(src_ack_net_1), .Y(
        src_ack_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hE) )  in_en_RNICUKI (.A(b6_nfs_IF[1]), .B(
        in_en_net_1), .Y(in_en_RNICUKI_net_1));
    CFG2 #( .INIT(4'h2) )  dout4_0_a2 (.A(dst_req_net_1), .B(
        dst_req_d_net_1), .Y(dout4));
    SLE \int_data[3]  (.D(b13_nAzGfFM_sLsv3_3), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[3]_net_1 ));
    CFG2 #( .INIT(4'hE) )  dout4_0_a2_RNIKLH5 (.A(b6_nfs_IF[1]), .B(
        dout4), .Y(dout4_0_a2_RNIKLH5_net_1));
    SLE src_req (.D(src_ack_i_0), .CLK(BW_clk_c), .EN(
        src_req_RNO_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        src_req_net_1));
    SLE dst_req_d (.D(dst_req_d_0), .CLK(IICE_comm2iice[11]), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dst_req_d_net_1));
    CFG2 #( .INIT(4'h4) )  dst_req_d_r (.A(b6_nfs_IF[1]), .B(
        dst_req_net_1), .Y(dst_req_d_0));
    
endmodule


module b7_OCByLXC_Z1_x_0(
       b6_Ocm0rW_0_0_o2,
       IICE_comm2iice,
       b13_nAzGfFM_sLsv3_0,
       b8_SoWGfWYY,
       b8_SoWGfWYY_i,
       BW_clk_c,
       b12_uRrc2XfY_Lyh,
       b11_PSyil9s_FMZ,
       b11_uRrc2XfY_XH,
       b4_PLyF,
       b13_nUTQBgfDb_Z4D,
       b12_nUTQBgfDb_bd,
       b16_nYhI39swMeEd_A78,
       b15_nYhI39swMeEd_Mg,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_XH
    );
output [2:2] b6_Ocm0rW_0_0_o2;
input  [11:8] IICE_comm2iice;
output b13_nAzGfFM_sLsv3_0;
output b8_SoWGfWYY;
output b8_SoWGfWYY_i;
input  BW_clk_c;
output b12_uRrc2XfY_Lyh;
input  b11_PSyil9s_FMZ;
input  b11_uRrc2XfY_XH;
input  b4_PLyF;
output b13_nUTQBgfDb_Z4D;
input  b12_nUTQBgfDb_bd;
output b16_nYhI39swMeEd_A78;
input  b15_nYhI39swMeEd_Mg;
output b12_vABZ3qsY_Lyh;
input  b11_vABZ3qsY_XH;

    wire \b13_nAzGfFM_sLsv3_i[0]_net_1 , \b13_nAzGfFM_sLsv3_i_i_0[0] , 
        \b3_nfs[0]_net_1 , VCC_net_1, \b6_nfs_IF[0] , GND_net_1, 
        \b3_nfs[1]_net_1 , \b6_nfs_IF[1] , \b3_nfs[2]_net_1 , 
        \b6_nfs_IF[2] , \b3_nfs[3]_net_1 , \b6_nfs_IF[3] , 
        \b3_nfs[4]_net_1 , \b6_nfs_IF[4] , 
        \b12_uRrc2XfY_rbN[19]_net_1 , \b12_uRrc2XfY_rbN_5[19]_net_1 , 
        un1_b12_uRrc2XfY_rbN10_i_0, \b12_uRrc2XfY_rbN[20]_net_1 , 
        \b12_uRrc2XfY_rbN_5[20]_net_1 , \b12_uRrc2XfY_rbN[21]_net_1 , 
        \b12_uRrc2XfY_rbN_5[21]_net_1 , \b12_uRrc2XfY_rbN[22]_net_1 , 
        \b12_uRrc2XfY_rbN_5[22]_net_1 , \b12_uRrc2XfY_rbN[23]_net_1 , 
        \b12_uRrc2XfY_rbN_5[23]_net_1 , \b12_uRrc2XfY_rbN[24]_net_1 , 
        \b12_uRrc2XfY_rbN_5[24]_net_1 , \b12_uRrc2XfY_rbN[25]_net_1 , 
        \b12_uRrc2XfY_rbN_5[25]_net_1 , \b12_uRrc2XfY_rbN[4]_net_1 , 
        \b12_uRrc2XfY_rbN_5[4]_net_1 , \b12_uRrc2XfY_rbN[5]_net_1 , 
        \b12_uRrc2XfY_rbN_5[5]_net_1 , \b12_uRrc2XfY_rbN[6]_net_1 , 
        \b12_uRrc2XfY_rbN_5[6]_net_1 , \b12_uRrc2XfY_rbN[7]_net_1 , 
        \b12_uRrc2XfY_rbN_5[7]_net_1 , \b12_uRrc2XfY_rbN[8]_net_1 , 
        \b12_uRrc2XfY_rbN_5[8]_net_1 , \b12_uRrc2XfY_rbN[9]_net_1 , 
        \b12_uRrc2XfY_rbN_5[9]_net_1 , \b12_uRrc2XfY_rbN[10]_net_1 , 
        \b12_uRrc2XfY_rbN_5[10]_net_1 , \b12_uRrc2XfY_rbN[11]_net_1 , 
        \b12_uRrc2XfY_rbN_5[11]_net_1 , \b12_uRrc2XfY_rbN[12]_net_1 , 
        \b12_uRrc2XfY_rbN_5[12]_net_1 , \b12_uRrc2XfY_rbN[13]_net_1 , 
        \b12_uRrc2XfY_rbN_5[13]_net_1 , \b12_uRrc2XfY_rbN[14]_net_1 , 
        \b12_uRrc2XfY_rbN_5[14]_net_1 , \b12_uRrc2XfY_rbN[15]_net_1 , 
        \b12_uRrc2XfY_rbN_5[15]_net_1 , \b12_uRrc2XfY_rbN[16]_net_1 , 
        \b12_uRrc2XfY_rbN_5[16]_net_1 , \b12_uRrc2XfY_rbN[17]_net_1 , 
        \b12_uRrc2XfY_rbN_5[17]_net_1 , \b12_uRrc2XfY_rbN[18]_net_1 , 
        \b12_uRrc2XfY_rbN_5[18]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[15]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[15]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[16]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[16]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[17]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[17]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[18]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[18]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[19]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[19]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[20]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[20]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[21]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[21]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[22]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[22]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[23]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[23]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[24]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[24]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[25]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[25]_net_1 , \b12_uRrc2XfY_rbN_5[0]_net_1 , 
        \b12_uRrc2XfY_rbN[1]_net_1 , \b12_uRrc2XfY_rbN_5[1]_net_1 , 
        \b12_uRrc2XfY_rbN[2]_net_1 , \b12_uRrc2XfY_rbN_5[2]_net_1 , 
        \b12_uRrc2XfY_rbN[3]_net_1 , \b12_uRrc2XfY_rbN_5[3]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[0]_net_1 , \b15_uRrc2XfY_rbN_gr[0]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[1]_net_1 , \b15_uRrc2XfY_rbN_gr[1]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[2]_net_1 , \b15_uRrc2XfY_rbN_gr[2]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[3]_net_1 , \b15_uRrc2XfY_rbN_gr[3]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[5]_net_1 , \b15_uRrc2XfY_rbN_gr[5]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[6]_net_1 , \b15_uRrc2XfY_rbN_gr[6]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[7]_net_1 , \b15_uRrc2XfY_rbN_gr[7]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[8]_net_1 , \b15_uRrc2XfY_rbN_gr[8]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[9]_net_1 , \b15_uRrc2XfY_rbN_gr[9]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[10]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[10]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[11]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[11]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[12]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[12]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[13]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[13]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[14]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[14]_net_1 , N_103_i_0, N_104_i_0, 
        \b13_nAzGfFM_sLsv3[5]_net_1 , b11_vABZ3qsY_qH, 
        \b7_nYhI39s[0]_net_1 , \b7_nYhI39s[1]_net_1 , 
        \b7_nYhI39s[2]_net_1 , \b7_nYhI39s[3]_net_1 , 
        \b7_nYhI39s[4]_net_1 , \b7_nYhI39s[5]_net_1 , 
        \b7_nYhI39s[6]_net_1 , \b7_nYhI39s[7]_net_1 , 
        \b7_nYhI39s[8]_net_1 , \b7_nYhI39s[9]_net_1 , 
        \status_b2sclk[0] , \status_b2sclk[1] , \status_b2sclk[2] , 
        \status_b2sclk[3] , \b13_nAzGfFM_sLsv3[2]_net_1 , 
        \b6_nfs_IF_i_0[1] , N_94_i_0, N_16, 
        \b13_nAzGfFM_sLsv3[3]_net_1 , N_90_i_0, 
        \b13_nAzGfFM_sLsv3[4]_net_1 , N_26_i_0, N_28_i_0, 
        b10_nYhI3_umjB_net_1, b10_nYhI3_umjB_3, 
        un1_b13_nAzGfFM_sLsv3_1_i_0, b8_vABZ3qsY_net_1, 
        \b3_nUT[8]_net_1 , \b6_nUT_IF[8] , \b3_nUT[9]_net_1 , 
        \b6_nUT_IF[9] , \b3_nUT[0]_net_1 , \b6_nUT_IF[0] , 
        \b3_nUT[1]_net_1 , \b6_nUT_IF[1] , \b3_nUT[2]_net_1 , 
        \b6_nUT_IF[2] , \b3_nUT[3]_net_1 , \b6_nUT_IF[3] , 
        \b3_nUT[4]_net_1 , \b6_nUT_IF[4] , \b3_nUT[5]_net_1 , 
        \b6_nUT_IF[5] , \b3_nUT[6]_net_1 , \b6_nUT_IF[6] , 
        \b3_nUT[7]_net_1 , \b6_nUT_IF[7] , \b7_nYhI39s_s[0] , N_23_i_0, 
        \b7_nYhI39s_s[1] , \b7_nYhI39s_s[2] , \b7_nYhI39s_s[3] , 
        \b7_nYhI39s_s[4] , \b7_nYhI39s_s[5] , \b7_nYhI39s_s[6] , 
        \b7_nYhI39s_s[7] , \b7_nYhI39s_s[8] , \b7_nYhI39s_s[9] , 
        b7_nYhI39s_cry_cy, \b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] , N_38, 
        \b7_nYhI39s_cry[0] , \b7_nYhI39s_5[0]_net_1 , 
        \b7_nYhI39s_cry[1] , \b7_nYhI39s_5[1]_net_1 , 
        \b7_nYhI39s_cry[2] , \b7_nYhI39s_5[2]_net_1 , 
        \b7_nYhI39s_cry[3] , \b7_nYhI39s_5[3]_net_1 , 
        \b7_nYhI39s_cry[4] , \b7_nYhI39s_5[4]_net_1 , 
        \b7_nYhI39s_cry[5] , \b7_nYhI39s_5[5]_net_1 , 
        \b7_nYhI39s_cry[6] , \b7_nYhI39s_5[6]_net_1 , 
        \b7_nYhI39s_cry[7] , \b7_nYhI39s_5[7]_net_1 , 
        \b7_nYhI39s_5[9]_net_1 , \b7_nYhI39s_cry[8] , 
        \b7_nYhI39s_5[8]_net_1 , 
        \b13_nAzGfFM_sLsv3_srsts_i_i_a2_0[2]_net_1 , G_60_4, 
        \b13_nAzGfFM_sLsv3_srsts_i_i_o2[2]_net_1 , G_60_6, G_60_5, 
        \b3_nfs_RNIPR5A1[2]_net_1 , 
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2[3]_net_1 , 
        \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]_net_1 , 
        \b6_Ocm0rW_0_i_a2_1[1]_net_1 , 
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]_net_1 , \b6_Ocm0rW[2] ;
    
    SLE \b3_nUT[0]  (.D(\b6_nUT_IF[0] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  b12_voSc3_gmasbb_RNO (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .Y(
        \b13_nAzGfFM_sLsv3_i_i_0[0] ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[2]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[2]_net_1 ), .Y(\b7_nYhI39s_5[2]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[6]  (.A(
        \b12_uRrc2XfY_rbN[7]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[6]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[6]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[12]  (.D(\b15_uRrc2XfY_rbN_gr[12]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[12]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[11]  (.D(\b12_uRrc2XfY_rbN_5[11]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[11]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[0]  (.D(\status_b2sclk[0] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[0]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  \b13_nAzGfFM_sLsv3_srsts_i_i_a2_0[2]  (
        .A(\b13_nAzGfFM_sLsv3[2]_net_1 ), .B(\b6_nfs_IF[1] ), .C(
        \b3_nfs[4]_net_1 ), .D(b11_PSyil9s_FMZ), .Y(
        \b13_nAzGfFM_sLsv3_srsts_i_i_a2_0[2]_net_1 ));
    b8_nR_ymqrG_10s_5s_0_0s_0s_1_510_x_0 b11_nUTGT_khWqH (
        .b6_nfs_IF_i_0({\b6_nfs_IF_i_0[1] }), .b6_nUT_IF({
        \b6_nUT_IF[9] , \b6_nUT_IF[8] , \b6_nUT_IF[7] , \b6_nUT_IF[6] , 
        \b6_nUT_IF[5] , \b6_nUT_IF[4] , \b6_nUT_IF[3] , \b6_nUT_IF[2] , 
        \b6_nUT_IF[1] , \b6_nUT_IF[0] }), .b6_nfs_IF({\b6_nfs_IF[4] , 
        \b6_nfs_IF[3] , \b6_nfs_IF[2] , \b6_nfs_IF[1] , \b6_nfs_IF[0] })
        , .IICE_comm2iice_3(IICE_comm2iice[11]), .IICE_comm2iice_0(
        IICE_comm2iice[8]), .IICE_comm2iice_2(IICE_comm2iice[10]), 
        .b4_PLyF(b4_PLyF), .b13_nUTQBgfDb_Z4D(b13_nUTQBgfDb_Z4D), 
        .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), .b16_nYhI39swMeEd_A78(
        b16_nYhI39swMeEd_A78), .b15_nYhI39swMeEd_Mg(
        b15_nYhI39swMeEd_Mg), .b12_vABZ3qsY_Lyh(b12_vABZ3qsY_Lyh), 
        .b11_vABZ3qsY_qH(b11_vABZ3qsY_qH), .b11_vABZ3qsY_XH(
        b11_vABZ3qsY_XH));
    SLE \b3_nUT[6]  (.D(\b6_nUT_IF[6] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[6]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \b6_Ocm0rW_0_0_o2[2]  (.A(
        \b13_nAzGfFM_sLsv3[2]_net_1 ), .B(\b13_nAzGfFM_sLsv3[3]_net_1 )
        , .Y(b6_Ocm0rW_0_0_o2[2]));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[17]  (.A(
        \b12_uRrc2XfY_rbN[18]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[17]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[17]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[4]  (.D(\b12_uRrc2XfY_rbN_5[4]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[4]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[0]  (.D(\b12_uRrc2XfY_rbN_5[0]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(b12_uRrc2XfY_Lyh));
    SLE \b15_uRrc2XfY_rbN_gs[1]  (.D(\b15_uRrc2XfY_rbN_gr[1]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[10]  (.D(\b15_uRrc2XfY_rbN_gr[10]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[10]_net_1 ));
    SLE \b3_nfs[1]  (.D(\b6_nfs_IF[1] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[5]  (.D(\b15_uRrc2XfY_rbN_gr[5]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \b6_Ocm0rW_0_0[2]  (.A(
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]_net_1 ), .B(
        b13_nAzGfFM_sLsv3_0), .C(b6_Ocm0rW_0_0_o2[2]), .Y(
        \b6_Ocm0rW[2] ));
    SLE \b15_uRrc2XfY_rbN_gr[18]  (.D(\b7_nYhI39s[2]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[18]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[14]  (.D(\b12_uRrc2XfY_rbN_5[14]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[14]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIF3AKE[3]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[3]_net_1 ), .D(\b7_nYhI39s_5[3]_net_1 ), .FCI(
        \b7_nYhI39s_cry[2] ), .S(\b7_nYhI39s_s[3] ), .Y(), .FCO(
        \b7_nYhI39s_cry[3] ));
    SLE \b7_nYhI39s[3]  (.D(\b7_nYhI39s_s[3] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[23]  (.D(\b7_nYhI39s[7]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[23]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[24]  (.D(\b15_uRrc2XfY_rbN_gr[24]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[24]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[13]  (.D(\b12_uRrc2XfY_rbN_5[13]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[13]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[1]  (.D(N_94_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b13_nAzGfFM_sLsv3_0));
    SLE \b12_uRrc2XfY_rbN[25]  (.D(\b12_uRrc2XfY_rbN_5[25]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[25]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[13]  (.D(N_104_i_0), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[13]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \b13_nAzGfFM_sLsv3_srsts_i_i_o2[2]  (.A(
        \b13_nAzGfFM_sLsv3[2]_net_1 ), .B(b11_PSyil9s_FMZ), .Y(
        \b13_nAzGfFM_sLsv3_srsts_i_i_o2[2]_net_1 ));
    CFG4 #( .INIT(16'hF0F8) )  \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]  (.A(
        \b13_nAzGfFM_sLsv3[2]_net_1 ), .B(b13_nAzGfFM_sLsv3_0), .C(
        \b13_nAzGfFM_sLsv3_srsts_i_i_a2_0[2]_net_1 ), .D(
        \b6_nfs_IF[1] ), .Y(\b13_nAzGfFM_sLsv3_srsts_i_i_0[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[19]  (.D(\b15_uRrc2XfY_rbN_gr[19]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[19]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[23]  (.A(
        \b12_uRrc2XfY_rbN[24]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[23]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[23]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[19]  (.D(\b12_uRrc2XfY_rbN_5[19]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[19]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[24]  (.A(
        \b12_uRrc2XfY_rbN[25]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[24]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[24]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[25]  (.D(\b15_uRrc2XfY_rbN_gr[25]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[25]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[6]  (.D(\b12_uRrc2XfY_rbN_5[6]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[6]_net_1 ));
    SLE \b3_nUT[1]  (.D(\b6_nUT_IF[1] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[17]  (.D(\b15_uRrc2XfY_rbN_gr[17]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[17]_net_1 ));
    CFG4 #( .INIT(16'h0A0E) )  \b13_nAzGfFM_sLsv3_RNO[4]  (.A(
        \b13_nAzGfFM_sLsv3[4]_net_1 ), .B(b10_nYhI3_umjB_net_1), .C(
        \b6_nfs_IF[1] ), .D(\b13_nAzGfFM_sLsv3_srsts_i_0_a2[3]_net_1 ), 
        .Y(N_26_i_0));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNI7BTMQ[7]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[7]_net_1 ), .D(\b7_nYhI39s_5[7]_net_1 ), .FCI(
        \b7_nYhI39s_cry[6] ), .S(\b7_nYhI39s_s[7] ), .Y(), .FCO(
        \b7_nYhI39s_cry[7] ));
    SLE \b7_nYhI39s[6]  (.D(\b7_nYhI39s_s[6] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[6]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[6]  (.D(\b15_uRrc2XfY_rbN_gr[6]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[6]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[14]  (.D(\b15_uRrc2XfY_rbN_gr[14]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[14]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[8]  (.D(\b12_uRrc2XfY_rbN_5[8]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[8]_net_1 ));
    CFG3 #( .INIT(8'hC8) )  un1_b12_uRrc2XfY_rbN10_i (.A(
        IICE_comm2iice[9]), .B(b11_uRrc2XfY_XH), .C(IICE_comm2iice[10])
        , .Y(un1_b12_uRrc2XfY_rbN10_i_0));
    SLE \b7_nYhI39s[5]  (.D(\b7_nYhI39s_s[5] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[5]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[1]  (.D(\b12_uRrc2XfY_rbN_5[1]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[3]  (.D(\status_b2sclk[3] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[3]_net_1 ));
    SLE \b3_nUT[3]  (.D(\b6_nUT_IF[3] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[15]  (.D(\b15_uRrc2XfY_rbN_gr[15]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[15]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[22]  (.D(\b7_nYhI39s[6]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[22]_net_1 ));
    CFG3 #( .INIT(8'hDF) )  b10_nYhI3_umjB_RNO_0 (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .B(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .C(N_38), .Y(
        un1_b13_nAzGfFM_sLsv3_1_i_0));
    SLE \b3_nfs[0]  (.D(\b6_nfs_IF[0] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[0]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[22]  (.A(
        \b12_uRrc2XfY_rbN[23]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[22]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[22]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[1]  (.A(
        \b12_uRrc2XfY_rbN[2]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[1]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[1]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3_i[0]  (.D(\b6_nfs_IF_i_0[1] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \b15_uRrc2XfY_rbN_gr_RNO[11]  (.A(
        \b13_nAzGfFM_sLsv3[5]_net_1 ), .B(\b13_nAzGfFM_sLsv3[3]_net_1 )
        , .C(b13_nAzGfFM_sLsv3_0), .Y(N_103_i_0));
    CFG4 #( .INIT(16'h0100) )  b10_nYhI3_umjB_RNO_3 (.A(
        \b7_nYhI39s[9]_net_1 ), .B(\b7_nYhI39s[6]_net_1 ), .C(
        \b7_nYhI39s[5]_net_1 ), .D(\b7_nYhI39s[0]_net_1 ), .Y(G_60_5));
    CFG2 #( .INIT(4'h1) )  b10_nYhI3_umjB_RNO_1 (.A(
        \b7_nYhI39s[3]_net_1 ), .B(\b7_nYhI39s[7]_net_1 ), .Y(G_60_4));
    SLE \b15_uRrc2XfY_rbN_gr[12]  (.D(b6_Ocm0rW_0_0_o2[2]), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[12]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[2]  (.A(
        \b12_uRrc2XfY_rbN[3]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[2]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[9]  (.D(\b15_uRrc2XfY_rbN_gr[9]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[9]_net_1 ));
    SLE \b7_nYhI39s[4]  (.D(\b7_nYhI39s_s[4] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[4]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[8]  (.A(
        \b12_uRrc2XfY_rbN[9]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[8]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[8]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[20]  (.D(\b7_nYhI39s[4]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[20]_net_1 ));
    ARI1 #( .INIT(20'h40E00) )  \b13_nAzGfFM_sLsv3_RNINSNH2[3]  (.A(
        VCC_net_1), .B(N_38), .C(b10_nYhI3_umjB_net_1), .D(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .FCI(VCC_net_1), .S(), .Y(
        \b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .FCO(b7_nYhI39s_cry_cy));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[5]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[5]_net_1 ), .Y(\b7_nYhI39s_5[5]_net_1 ));
    SLE \b7_nYhI39s[9]  (.D(\b7_nYhI39s_s[9] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[9]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \b3_nfs_RNIPR5A1[2]  (.A(\b3_nfs[2]_net_1 )
        , .B(\b3_nfs[4]_net_1 ), .C(\b3_nfs[3]_net_1 ), .Y(
        \b3_nfs_RNIPR5A1[2]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[15]  (.D(\b12_uRrc2XfY_rbN_5[15]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[15]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[11]  (.A(
        \b12_uRrc2XfY_rbN[12]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[11]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[11]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \b13_nAzGfFM_sLsv3_RNO[5]  (.A(
        \b13_nAzGfFM_sLsv3[5]_net_1 ), .B(\b3_nfs[4]_net_1 ), .C(
        \b13_nAzGfFM_sLsv3_srsts_i_i_o2[2]_net_1 ), .D(\b6_nfs_IF[1] ), 
        .Y(N_28_i_0));
    SLE \b15_uRrc2XfY_rbN_gr[10]  (.D(\b6_nfs_IF[4] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[10]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]  (.A(
        b8_vABZ3qsY_net_1), .B(\b3_nfs[0]_net_1 ), .C(
        \b6_Ocm0rW_0_i_a2_1[1]_net_1 ), .Y(
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]_net_1 ));
    CFG3 #( .INIT(8'h07) )  \b13_nAzGfFM_sLsv3_srsts_i_0_a2[3]  (.A(
        b11_PSyil9s_FMZ), .B(\b13_nAzGfFM_sLsv3[2]_net_1 ), .C(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .Y(
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2[3]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNI7JJLK[5]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[5]_net_1 ), .D(\b7_nYhI39s_5[5]_net_1 ), .FCI(
        \b7_nYhI39s_cry[4] ), .S(\b7_nYhI39s_s[5] ), .Y(), .FCO(
        \b7_nYhI39s_cry[5] ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[15]  (.A(
        \b12_uRrc2XfY_rbN[16]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[15]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[15]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[10]  (.A(
        \b12_uRrc2XfY_rbN[11]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[10]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[10]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[0]  (.A(
        \b12_uRrc2XfY_rbN[1]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[0]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[0]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[6]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[6]_net_1 ), .Y(\b7_nYhI39s_5[6]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[5]  (.D(N_28_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[5]_net_1 ));
    CFG4 #( .INIT(16'h5FDF) )  b8_vABZ3qsY_RNIG4T32 (.A(
        b13_nAzGfFM_sLsv3_0), .B(\b3_nfs_RNIPR5A1[2]_net_1 ), .C(
        b8_vABZ3qsY_net_1), .D(\b3_nfs[0]_net_1 ), .Y(N_38));
    SLE \b15_uRrc2XfY_rbN_gs[21]  (.D(\b15_uRrc2XfY_rbN_gr[21]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[21]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[0]  (.D(\b15_uRrc2XfY_rbN_gr[0]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[0]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[18]  (.A(
        \b12_uRrc2XfY_rbN[19]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[18]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[18]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[7]  (.D(\b6_nfs_IF[1] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[8]  (.D(\b15_uRrc2XfY_rbN_gr[8]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[8]_net_1 ));
    clock2_en_reg_en_5s_x_0 iclksync (.IICE_comm2iice({
        IICE_comm2iice[11]}), .b6_nfs_IF_i_0({\b6_nfs_IF_i_0[1] }), 
        .status_b2sclk({\status_b2sclk[3] , \status_b2sclk[2] , 
        \status_b2sclk[1] , \status_b2sclk[0] }), .b6_nfs_IF({
        \b6_nfs_IF[1] }), .b6_Ocm0rW({\b6_Ocm0rW[2] }), 
        .b6_Ocm0rW_0_i_a2_1({\b6_Ocm0rW_0_i_a2_1[1]_net_1 }), 
        .b13_nAzGfFM_sLsv3_3(\b13_nAzGfFM_sLsv3[5]_net_1 ), 
        .b13_nAzGfFM_sLsv3_0(\b13_nAzGfFM_sLsv3[2]_net_1 ), 
        .b13_nAzGfFM_sLsv3_2(\b13_nAzGfFM_sLsv3[4]_net_1 ), .BW_clk_c(
        BW_clk_c), .N_38(N_38));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIAAINT[8]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[8]_net_1 ), .D(\b7_nYhI39s_5[8]_net_1 ), .FCI(
        \b7_nYhI39s_cry[7] ), .S(\b7_nYhI39s_s[8] ), .Y(), .FCO(
        \b7_nYhI39s_cry[8] ));
    SLE b12_voSc3_gmasbb (.D(\b13_nAzGfFM_sLsv3_i_i_0[0] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b8_SoWGfWYY));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[7]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[7]_net_1 ), .Y(\b7_nYhI39s_5[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[6]  (.D(\b6_nfs_IF[0] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[6]_net_1 ));
    SLE \b3_nUT[9]  (.D(\b6_nUT_IF[9] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[9]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[19]  (.D(\b7_nYhI39s[3]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[19]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \b6_Ocm0rW_0_i_a2_1[1]  (.A(
        b10_nYhI3_umjB_net_1), .B(\b3_nfs_RNIPR5A1[2]_net_1 ), .C(
        \b3_nfs[1]_net_1 ), .Y(\b6_Ocm0rW_0_i_a2_1[1]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[8]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[8]_net_1 ), .Y(\b7_nYhI39s_5[8]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[4]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[4]_net_1 ), .Y(\b7_nYhI39s_5[4]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[24]  (.D(\b7_nYhI39s[8]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[24]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[9]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[9]_net_1 ), .Y(\b7_nYhI39s_5[9]_net_1 ));
    SLE \b7_nYhI39s[0]  (.D(\b7_nYhI39s_s[0] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[0]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[5]  (.D(\b12_uRrc2XfY_rbN_5[5]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[5]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[18]  (.D(\b12_uRrc2XfY_rbN_5[18]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[18]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[16]  (.D(\b15_uRrc2XfY_rbN_gr[16]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[16]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[7]  (.A(
        \b12_uRrc2XfY_rbN[8]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[7]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[7]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[3]  (.D(\b12_uRrc2XfY_rbN_5[3]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[17]  (.D(\b7_nYhI39s[1]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[17]_net_1 ));
    SLE \b7_nYhI39s[2]  (.D(\b7_nYhI39s_s[2] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[2]  (.D(\b15_uRrc2XfY_rbN_gr[2]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[2]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \b15_uRrc2XfY_rbN_gr_RNO[13]  (.A(
        \b13_nAzGfFM_sLsv3[4]_net_1 ), .B(\b13_nAzGfFM_sLsv3[5]_net_1 )
        , .Y(N_104_i_0));
    SLE \b7_nYhI39s[8]  (.D(\b7_nYhI39s_s[8] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[8]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[11]  (.D(\b15_uRrc2XfY_rbN_gr[11]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[11]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[14]  (.D(\b13_nAzGfFM_sLsv3[5]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gr[14]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[3]  (.D(\b15_uRrc2XfY_rbN_gr[3]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[3]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[3]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[3]_net_1 ), .Y(\b7_nYhI39s_5[3]_net_1 ));
    SLE \b3_nUT[5]  (.D(\b6_nUT_IF[5] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[5]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  b10_nYhI3_umjB_RNO (.A(G_60_4), .B(
        G_60_6), .C(G_60_5), .D(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .Y(
        b10_nYhI3_umjB_3));
    SLE \b12_uRrc2XfY_rbN[22]  (.D(\b12_uRrc2XfY_rbN_5[22]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[22]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \b13_nAzGfFM_sLsv3_RNO[3]  (.A(
        b10_nYhI3_umjB_net_1), .B(\b6_nfs_IF[1] ), .C(
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2[3]_net_1 ), .Y(N_90_i_0));
    SLE \b3_nfs[4]  (.D(\b6_nfs_IF[4] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[4]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[8]  (.D(\b6_nfs_IF[2] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[8]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[3]  (.A(
        \b12_uRrc2XfY_rbN[4]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[3]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[3]_net_1 ));
    SLE \b3_nfs[2]  (.D(\b6_nfs_IF[2] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[25]  (.D(\b7_nYhI39s[9]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[25]_net_1 ));
    SLE \b3_nUT[8]  (.D(\b6_nUT_IF[8] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[8]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[20]  (.D(\b12_uRrc2XfY_rbN_5[20]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[20]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[9]  (.D(\b12_uRrc2XfY_rbN_5[9]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[9]_net_1 ));
    CFG1 #( .INIT(2'h1) )  b12_voSc3_gmasbb_RNIALH6 (.A(b8_SoWGfWYY), 
        .Y(b8_SoWGfWYY_i));
    SLE \b15_uRrc2XfY_rbN_gs[23]  (.D(\b15_uRrc2XfY_rbN_gr[23]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[23]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[16]  (.A(
        \b12_uRrc2XfY_rbN[17]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[16]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[16]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[15]  (.D(b11_vABZ3qsY_qH), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[15]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[4]  (.D(N_26_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[4]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[2]  (.D(\b12_uRrc2XfY_rbN_5[2]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[2]_net_1 ));
    CFG4 #( .INIT(16'h1311) )  \b13_nAzGfFM_sLsv3_RNO[1]  (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .B(\b6_nfs_IF[1] ), .C(
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]_net_1 ), .D(
        b13_nAzGfFM_sLsv3_0), .Y(N_94_i_0));
    SLE \b3_nUT[7]  (.D(\b6_nUT_IF[7] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[18]  (.D(\b15_uRrc2XfY_rbN_gr[18]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[18]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[19]  (.A(
        \b12_uRrc2XfY_rbN[20]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[19]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[19]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[21]  (.D(\b12_uRrc2XfY_rbN_5[21]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[21]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[13]  (.A(
        \b12_uRrc2XfY_rbN[14]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[13]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[13]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[14]  (.A(
        \b12_uRrc2XfY_rbN[15]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[14]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[14]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIABCI5[0]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[0]_net_1 ), .D(\b7_nYhI39s_5[0]_net_1 ), .FCI(
        b7_nYhI39s_cry_cy), .S(\b7_nYhI39s_s[0] ), .Y(), .FCO(
        \b7_nYhI39s_cry[0] ));
    SLE \b15_uRrc2XfY_rbN_gs[13]  (.D(\b15_uRrc2XfY_rbN_gr[13]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[13]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  b10_nYhI3_umjB_RNO_2 (.A(
        \b7_nYhI39s[8]_net_1 ), .B(\b7_nYhI39s[4]_net_1 ), .C(
        \b7_nYhI39s[2]_net_1 ), .D(\b7_nYhI39s[1]_net_1 ), .Y(G_60_6));
    CFG4 #( .INIT(16'h1D3F) )  \b13_nAzGfFM_sLsv3_i_RNIST5R2[0]  (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .B(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .C(b10_nYhI3_umjB_net_1), .D(
        N_38), .Y(N_23_i_0));
    SLE \b12_uRrc2XfY_rbN[16]  (.D(\b12_uRrc2XfY_rbN_5[16]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[16]_net_1 ));
    SLE b10_nYhI3_umjB (.D(b10_nYhI3_umjB_3), .CLK(BW_clk_c), .EN(
        un1_b13_nAzGfFM_sLsv3_1_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b10_nYhI3_umjB_net_1));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[0]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[0]_net_1 ), .Y(\b7_nYhI39s_5[0]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[1]  (.D(\status_b2sclk[1] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[1]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[5]  (.A(
        \b12_uRrc2XfY_rbN[6]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[5]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[5]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIAQUKH[4]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[4]_net_1 ), .D(\b7_nYhI39s_5[4]_net_1 ), .FCI(
        \b7_nYhI39s_cry[3] ), .S(\b7_nYhI39s_s[4] ), .Y(), .FCO(
        \b7_nYhI39s_cry[4] ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIMELJB[2]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[2]_net_1 ), .D(\b7_nYhI39s_5[2]_net_1 ), .FCI(
        \b7_nYhI39s_cry[1] ), .S(\b7_nYhI39s_s[2] ), .Y(), .FCO(
        \b7_nYhI39s_cry[2] ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIVR0J8[1]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[1]_net_1 ), .D(\b7_nYhI39s_5[1]_net_1 ), .FCI(
        \b7_nYhI39s_cry[0] ), .S(\b7_nYhI39s_s[1] ), .Y(), .FCO(
        \b7_nYhI39s_cry[1] ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[21]  (.A(
        \b12_uRrc2XfY_rbN[22]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[21]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[21]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[17]  (.D(\b12_uRrc2XfY_rbN_5[17]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[17]_net_1 ));
    SLE b8_vABZ3qsY (.D(b11_vABZ3qsY_qH), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b8_vABZ3qsY_net_1));
    SLE \b12_uRrc2XfY_rbN[24]  (.D(\b12_uRrc2XfY_rbN_5[24]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[24]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNI6E8MN[6]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[6]_net_1 ), .D(\b7_nYhI39s_5[6]_net_1 ), .FCI(
        \b7_nYhI39s_cry[5] ), .S(\b7_nYhI39s_s[6] ), .Y(), .FCO(
        \b7_nYhI39s_cry[6] ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[9]  (.A(
        \b12_uRrc2XfY_rbN[10]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[9]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[9]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[23]  (.D(\b12_uRrc2XfY_rbN_5[23]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[23]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[22]  (.D(\b15_uRrc2XfY_rbN_gr[22]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[22]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[12]  (.D(\b12_uRrc2XfY_rbN_5[12]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[12]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[2]  (.D(N_16), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[2]_net_1 ));
    ARI1 #( .INIT(20'h41B00) )  \b7_nYhI39s_RNO[9]  (.A(VCC_net_1), .B(
        \b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(\b7_nYhI39s[9]_net_1 ), 
        .D(\b7_nYhI39s_5[9]_net_1 ), .FCI(\b7_nYhI39s_cry[8] ), .S(
        \b7_nYhI39s_s[9] ), .Y(), .FCO());
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[25]  (.A(b4_PLyF), .B(
        IICE_comm2iice[9]), .C(\b15_uRrc2XfY_rbN_gs[25]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[25]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[20]  (.A(
        \b12_uRrc2XfY_rbN[21]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[20]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[20]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[12]  (.A(
        \b12_uRrc2XfY_rbN[13]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[12]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[12]_net_1 ));
    SLE \b3_nUT[2]  (.D(\b6_nUT_IF[2] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[2]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[10]  (.D(\b12_uRrc2XfY_rbN_5[10]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[10]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[9]  (.D(\b6_nfs_IF[3] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[9]_net_1 ));
    CFG3 #( .INIT(8'hFD) )  \b7_nYhI39s_5[1]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[1]_net_1 ), .Y(\b7_nYhI39s_5[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \b12_uRrc2XfY_rbN_5[4]  (.A(
        IICE_comm2iice[9]), .B(\b12_uRrc2XfY_rbN[5]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[4]_net_1 ));
    SLE \b3_nfs[3]  (.D(\b6_nfs_IF[3] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[21]  (.D(\b7_nYhI39s[5]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[21]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[7]  (.D(\b12_uRrc2XfY_rbN_5[7]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[7]_net_1 ));
    CFG4 #( .INIT(16'hAAEA) )  \b13_nAzGfFM_sLsv3_srsts_i_i[2]  (.A(
        \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]_net_1 ), .B(
        \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]_net_1 ), .C(
        b13_nAzGfFM_sLsv3_0), .D(\b6_nfs_IF[1] ), .Y(N_16));
    SLE \b13_nAzGfFM_sLsv3[3]  (.D(N_90_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[3]_net_1 ));
    SLE \b7_nYhI39s[1]  (.D(\b7_nYhI39s_s[1] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[20]  (.D(\b15_uRrc2XfY_rbN_gr[20]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[20]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[16]  (.D(\b7_nYhI39s[0]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[16]_net_1 ));
    SLE \b7_nYhI39s[7]  (.D(\b7_nYhI39s_s[7] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[7]  (.D(\b15_uRrc2XfY_rbN_gr[7]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[7]_net_1 ));
    SLE \b3_nUT[4]  (.D(\b6_nUT_IF[4] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[4]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[5]  (.D(\b13_nAzGfFM_sLsv3[2]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gr[5]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[2]  (.D(\status_b2sclk[2] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[11]  (.D(N_103_i_0), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[11]_net_1 ));
    
endmodule


module b3_12m_x_0(
       b6_Ocm0rW_0_0_o2,
       b13_nAzGfFM_sLsv3,
       IICE_comm2iice,
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b8_SoWGfWYY,
       b8_SoWGfWYY_i,
       BW_clk_c,
       b12_uRrc2XfY_Lyh,
       b11_PSyil9s_FMZ,
       b11_uRrc2XfY_XH,
       b4_PLyF,
       b13_nUTQBgfDb_Z4D,
       b12_nUTQBgfDb_bd,
       b16_nYhI39swMeEd_A78,
       b15_nYhI39swMeEd_Mg,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_XH,
       b7_PSyi3wy,
       b8_PSyiBgYG
    );
output [2:2] b6_Ocm0rW_0_0_o2;
output [1:1] b13_nAzGfFM_sLsv3;
input  [11:8] IICE_comm2iice;
input  [376:0] mdiclink_reg;
input  [376:0] b11_OFWNT9L_8tZ;
output b8_SoWGfWYY;
output b8_SoWGfWYY_i;
input  BW_clk_c;
output b12_uRrc2XfY_Lyh;
output b11_PSyil9s_FMZ;
input  b11_uRrc2XfY_XH;
input  b4_PLyF;
output b13_nUTQBgfDb_Z4D;
input  b12_nUTQBgfDb_bd;
output b16_nYhI39swMeEd_A78;
input  b15_nYhI39swMeEd_Mg;
output b12_vABZ3qsY_Lyh;
input  b11_vABZ3qsY_XH;
output b7_PSyi3wy;
input  b8_PSyiBgYG;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    b7_PfFzrNY_x_0 b4_PfFz (.mdiclink_reg({mdiclink_reg[376], 
        mdiclink_reg[375], mdiclink_reg[374], mdiclink_reg[373], 
        mdiclink_reg[372], mdiclink_reg[371], mdiclink_reg[370], 
        mdiclink_reg[369], mdiclink_reg[368], mdiclink_reg[367], 
        mdiclink_reg[366], mdiclink_reg[365], mdiclink_reg[364], 
        mdiclink_reg[363], mdiclink_reg[362], mdiclink_reg[361], 
        mdiclink_reg[360], mdiclink_reg[359], mdiclink_reg[358], 
        mdiclink_reg[357], mdiclink_reg[356], mdiclink_reg[355], 
        mdiclink_reg[354], mdiclink_reg[353], mdiclink_reg[352], 
        mdiclink_reg[351], mdiclink_reg[350], mdiclink_reg[349], 
        mdiclink_reg[348], mdiclink_reg[347], mdiclink_reg[346], 
        mdiclink_reg[345], mdiclink_reg[344], mdiclink_reg[343], 
        mdiclink_reg[342], mdiclink_reg[341], mdiclink_reg[340], 
        mdiclink_reg[339], mdiclink_reg[338], mdiclink_reg[337], 
        mdiclink_reg[336], mdiclink_reg[335], mdiclink_reg[334], 
        mdiclink_reg[333], mdiclink_reg[332], mdiclink_reg[331], 
        mdiclink_reg[330], mdiclink_reg[329], mdiclink_reg[328], 
        mdiclink_reg[327], mdiclink_reg[326], mdiclink_reg[325], 
        mdiclink_reg[324], mdiclink_reg[323], mdiclink_reg[322], 
        mdiclink_reg[321], mdiclink_reg[320], mdiclink_reg[319], 
        mdiclink_reg[318], mdiclink_reg[317], mdiclink_reg[316], 
        mdiclink_reg[315], mdiclink_reg[314], mdiclink_reg[313], 
        mdiclink_reg[312], mdiclink_reg[311], mdiclink_reg[310], 
        mdiclink_reg[309], mdiclink_reg[308], mdiclink_reg[307], 
        mdiclink_reg[306], mdiclink_reg[305], mdiclink_reg[304], 
        mdiclink_reg[303], mdiclink_reg[302], mdiclink_reg[301], 
        mdiclink_reg[300], mdiclink_reg[299], mdiclink_reg[298], 
        mdiclink_reg[297], mdiclink_reg[296], mdiclink_reg[295], 
        mdiclink_reg[294], mdiclink_reg[293], mdiclink_reg[292], 
        mdiclink_reg[291], mdiclink_reg[290], mdiclink_reg[289], 
        mdiclink_reg[288], mdiclink_reg[287], mdiclink_reg[286], 
        mdiclink_reg[285], mdiclink_reg[284], mdiclink_reg[283], 
        mdiclink_reg[282], mdiclink_reg[281], mdiclink_reg[280], 
        mdiclink_reg[279], mdiclink_reg[278], mdiclink_reg[277], 
        mdiclink_reg[276], mdiclink_reg[275], mdiclink_reg[274], 
        mdiclink_reg[273], mdiclink_reg[272], mdiclink_reg[271], 
        mdiclink_reg[270], mdiclink_reg[269], mdiclink_reg[268], 
        mdiclink_reg[267], mdiclink_reg[266], mdiclink_reg[265], 
        mdiclink_reg[264], mdiclink_reg[263], mdiclink_reg[262], 
        mdiclink_reg[261], mdiclink_reg[260], mdiclink_reg[259], 
        mdiclink_reg[258], mdiclink_reg[257], mdiclink_reg[256], 
        mdiclink_reg[255], mdiclink_reg[254], mdiclink_reg[253], 
        mdiclink_reg[252], mdiclink_reg[251], mdiclink_reg[250], 
        mdiclink_reg[249], mdiclink_reg[248], mdiclink_reg[247], 
        mdiclink_reg[246], mdiclink_reg[245], mdiclink_reg[244], 
        mdiclink_reg[243], mdiclink_reg[242], mdiclink_reg[241], 
        mdiclink_reg[240], mdiclink_reg[239], mdiclink_reg[238], 
        mdiclink_reg[237], mdiclink_reg[236], mdiclink_reg[235], 
        mdiclink_reg[234], mdiclink_reg[233], mdiclink_reg[232], 
        mdiclink_reg[231], mdiclink_reg[230], mdiclink_reg[229], 
        mdiclink_reg[228], mdiclink_reg[227], mdiclink_reg[226], 
        mdiclink_reg[225], mdiclink_reg[224], mdiclink_reg[223], 
        mdiclink_reg[222], mdiclink_reg[221], mdiclink_reg[220], 
        mdiclink_reg[219], mdiclink_reg[218], mdiclink_reg[217], 
        mdiclink_reg[216], mdiclink_reg[215], mdiclink_reg[214], 
        mdiclink_reg[213], mdiclink_reg[212], mdiclink_reg[211], 
        mdiclink_reg[210], mdiclink_reg[209], mdiclink_reg[208], 
        mdiclink_reg[207], mdiclink_reg[206], mdiclink_reg[205], 
        mdiclink_reg[204], mdiclink_reg[203], mdiclink_reg[202], 
        mdiclink_reg[201], mdiclink_reg[200], mdiclink_reg[199], 
        mdiclink_reg[198], mdiclink_reg[197], mdiclink_reg[196], 
        mdiclink_reg[195], mdiclink_reg[194], mdiclink_reg[193], 
        mdiclink_reg[192], mdiclink_reg[191], mdiclink_reg[190], 
        mdiclink_reg[189], mdiclink_reg[188], mdiclink_reg[187], 
        mdiclink_reg[186], mdiclink_reg[185], mdiclink_reg[184], 
        mdiclink_reg[183], mdiclink_reg[182], mdiclink_reg[181], 
        mdiclink_reg[180], mdiclink_reg[179], mdiclink_reg[178], 
        mdiclink_reg[177], mdiclink_reg[176], mdiclink_reg[175], 
        mdiclink_reg[174], mdiclink_reg[173], mdiclink_reg[172], 
        mdiclink_reg[171], mdiclink_reg[170], mdiclink_reg[169], 
        mdiclink_reg[168], mdiclink_reg[167], mdiclink_reg[166], 
        mdiclink_reg[165], mdiclink_reg[164], mdiclink_reg[163], 
        mdiclink_reg[162], mdiclink_reg[161], mdiclink_reg[160], 
        mdiclink_reg[159], mdiclink_reg[158], mdiclink_reg[157], 
        mdiclink_reg[156], mdiclink_reg[155], mdiclink_reg[154], 
        mdiclink_reg[153], mdiclink_reg[152], mdiclink_reg[151], 
        mdiclink_reg[150], mdiclink_reg[149], mdiclink_reg[148], 
        mdiclink_reg[147], mdiclink_reg[146], mdiclink_reg[145], 
        mdiclink_reg[144], mdiclink_reg[143], mdiclink_reg[142], 
        mdiclink_reg[141], mdiclink_reg[140], mdiclink_reg[139], 
        mdiclink_reg[138], mdiclink_reg[137], mdiclink_reg[136], 
        mdiclink_reg[135], mdiclink_reg[134], mdiclink_reg[133], 
        mdiclink_reg[132], mdiclink_reg[131], mdiclink_reg[130], 
        mdiclink_reg[129], mdiclink_reg[128], mdiclink_reg[127], 
        mdiclink_reg[126], mdiclink_reg[125], mdiclink_reg[124], 
        mdiclink_reg[123], mdiclink_reg[122], mdiclink_reg[121], 
        mdiclink_reg[120], mdiclink_reg[119], mdiclink_reg[118], 
        mdiclink_reg[117], mdiclink_reg[116], mdiclink_reg[115], 
        mdiclink_reg[114], mdiclink_reg[113], mdiclink_reg[112], 
        mdiclink_reg[111], mdiclink_reg[110], mdiclink_reg[109], 
        mdiclink_reg[108], mdiclink_reg[107], mdiclink_reg[106], 
        mdiclink_reg[105], mdiclink_reg[104], mdiclink_reg[103], 
        mdiclink_reg[102], mdiclink_reg[101], mdiclink_reg[100], 
        mdiclink_reg[99], mdiclink_reg[98], mdiclink_reg[97], 
        mdiclink_reg[96], mdiclink_reg[95], mdiclink_reg[94], 
        mdiclink_reg[93], mdiclink_reg[92], mdiclink_reg[91], 
        mdiclink_reg[90], mdiclink_reg[89], mdiclink_reg[88], 
        mdiclink_reg[87], mdiclink_reg[86], mdiclink_reg[85], 
        mdiclink_reg[84], mdiclink_reg[83], mdiclink_reg[82], 
        mdiclink_reg[81], mdiclink_reg[80], mdiclink_reg[79], 
        mdiclink_reg[78], mdiclink_reg[77], mdiclink_reg[76], 
        mdiclink_reg[75], mdiclink_reg[74], mdiclink_reg[73], 
        mdiclink_reg[72], mdiclink_reg[71], mdiclink_reg[70], 
        mdiclink_reg[69], mdiclink_reg[68], mdiclink_reg[67], 
        mdiclink_reg[66], mdiclink_reg[65], mdiclink_reg[64], 
        mdiclink_reg[63], mdiclink_reg[62], mdiclink_reg[61], 
        mdiclink_reg[60], mdiclink_reg[59], mdiclink_reg[58], 
        mdiclink_reg[57], mdiclink_reg[56], mdiclink_reg[55], 
        mdiclink_reg[54], mdiclink_reg[53], mdiclink_reg[52], 
        mdiclink_reg[51], mdiclink_reg[50], mdiclink_reg[49], 
        mdiclink_reg[48], mdiclink_reg[47], mdiclink_reg[46], 
        mdiclink_reg[45], mdiclink_reg[44], mdiclink_reg[43], 
        mdiclink_reg[42], mdiclink_reg[41], mdiclink_reg[40], 
        mdiclink_reg[39], mdiclink_reg[38], mdiclink_reg[37], 
        mdiclink_reg[36], mdiclink_reg[35], mdiclink_reg[34], 
        mdiclink_reg[33], mdiclink_reg[32], mdiclink_reg[31], 
        mdiclink_reg[30], mdiclink_reg[29], mdiclink_reg[28], 
        mdiclink_reg[27], mdiclink_reg[26], mdiclink_reg[25], 
        mdiclink_reg[24], mdiclink_reg[23], mdiclink_reg[22], 
        mdiclink_reg[21], mdiclink_reg[20], mdiclink_reg[19], 
        mdiclink_reg[18], mdiclink_reg[17], mdiclink_reg[16], 
        mdiclink_reg[15], mdiclink_reg[14], mdiclink_reg[13], 
        mdiclink_reg[12], mdiclink_reg[11], mdiclink_reg[10], 
        mdiclink_reg[9], mdiclink_reg[8], mdiclink_reg[7], 
        mdiclink_reg[6], mdiclink_reg[5], mdiclink_reg[4], 
        mdiclink_reg[3], mdiclink_reg[2], mdiclink_reg[1], 
        mdiclink_reg[0]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[376], 
        b11_OFWNT9L_8tZ[375], b11_OFWNT9L_8tZ[374], 
        b11_OFWNT9L_8tZ[373], b11_OFWNT9L_8tZ[372], 
        b11_OFWNT9L_8tZ[371], b11_OFWNT9L_8tZ[370], 
        b11_OFWNT9L_8tZ[369], b11_OFWNT9L_8tZ[368], 
        b11_OFWNT9L_8tZ[367], b11_OFWNT9L_8tZ[366], 
        b11_OFWNT9L_8tZ[365], b11_OFWNT9L_8tZ[364], 
        b11_OFWNT9L_8tZ[363], b11_OFWNT9L_8tZ[362], 
        b11_OFWNT9L_8tZ[361], b11_OFWNT9L_8tZ[360], 
        b11_OFWNT9L_8tZ[359], b11_OFWNT9L_8tZ[358], 
        b11_OFWNT9L_8tZ[357], b11_OFWNT9L_8tZ[356], 
        b11_OFWNT9L_8tZ[355], b11_OFWNT9L_8tZ[354], 
        b11_OFWNT9L_8tZ[353], b11_OFWNT9L_8tZ[352], 
        b11_OFWNT9L_8tZ[351], b11_OFWNT9L_8tZ[350], 
        b11_OFWNT9L_8tZ[349], b11_OFWNT9L_8tZ[348], 
        b11_OFWNT9L_8tZ[347], b11_OFWNT9L_8tZ[346], 
        b11_OFWNT9L_8tZ[345], b11_OFWNT9L_8tZ[344], 
        b11_OFWNT9L_8tZ[343], b11_OFWNT9L_8tZ[342], 
        b11_OFWNT9L_8tZ[341], b11_OFWNT9L_8tZ[340], 
        b11_OFWNT9L_8tZ[339], b11_OFWNT9L_8tZ[338], 
        b11_OFWNT9L_8tZ[337], b11_OFWNT9L_8tZ[336], 
        b11_OFWNT9L_8tZ[335], b11_OFWNT9L_8tZ[334], 
        b11_OFWNT9L_8tZ[333], b11_OFWNT9L_8tZ[332], 
        b11_OFWNT9L_8tZ[331], b11_OFWNT9L_8tZ[330], 
        b11_OFWNT9L_8tZ[329], b11_OFWNT9L_8tZ[328], 
        b11_OFWNT9L_8tZ[327], b11_OFWNT9L_8tZ[326], 
        b11_OFWNT9L_8tZ[325], b11_OFWNT9L_8tZ[324], 
        b11_OFWNT9L_8tZ[323], b11_OFWNT9L_8tZ[322], 
        b11_OFWNT9L_8tZ[321], b11_OFWNT9L_8tZ[320], 
        b11_OFWNT9L_8tZ[319], b11_OFWNT9L_8tZ[318], 
        b11_OFWNT9L_8tZ[317], b11_OFWNT9L_8tZ[316], 
        b11_OFWNT9L_8tZ[315], b11_OFWNT9L_8tZ[314], 
        b11_OFWNT9L_8tZ[313], b11_OFWNT9L_8tZ[312], 
        b11_OFWNT9L_8tZ[311], b11_OFWNT9L_8tZ[310], 
        b11_OFWNT9L_8tZ[309], b11_OFWNT9L_8tZ[308], 
        b11_OFWNT9L_8tZ[307], b11_OFWNT9L_8tZ[306], 
        b11_OFWNT9L_8tZ[305], b11_OFWNT9L_8tZ[304], 
        b11_OFWNT9L_8tZ[303], b11_OFWNT9L_8tZ[302], 
        b11_OFWNT9L_8tZ[301], b11_OFWNT9L_8tZ[300], 
        b11_OFWNT9L_8tZ[299], b11_OFWNT9L_8tZ[298], 
        b11_OFWNT9L_8tZ[297], b11_OFWNT9L_8tZ[296], 
        b11_OFWNT9L_8tZ[295], b11_OFWNT9L_8tZ[294], 
        b11_OFWNT9L_8tZ[293], b11_OFWNT9L_8tZ[292], 
        b11_OFWNT9L_8tZ[291], b11_OFWNT9L_8tZ[290], 
        b11_OFWNT9L_8tZ[289], b11_OFWNT9L_8tZ[288], 
        b11_OFWNT9L_8tZ[287], b11_OFWNT9L_8tZ[286], 
        b11_OFWNT9L_8tZ[285], b11_OFWNT9L_8tZ[284], 
        b11_OFWNT9L_8tZ[283], b11_OFWNT9L_8tZ[282], 
        b11_OFWNT9L_8tZ[281], b11_OFWNT9L_8tZ[280], 
        b11_OFWNT9L_8tZ[279], b11_OFWNT9L_8tZ[278], 
        b11_OFWNT9L_8tZ[277], b11_OFWNT9L_8tZ[276], 
        b11_OFWNT9L_8tZ[275], b11_OFWNT9L_8tZ[274], 
        b11_OFWNT9L_8tZ[273], b11_OFWNT9L_8tZ[272], 
        b11_OFWNT9L_8tZ[271], b11_OFWNT9L_8tZ[270], 
        b11_OFWNT9L_8tZ[269], b11_OFWNT9L_8tZ[268], 
        b11_OFWNT9L_8tZ[267], b11_OFWNT9L_8tZ[266], 
        b11_OFWNT9L_8tZ[265], b11_OFWNT9L_8tZ[264], 
        b11_OFWNT9L_8tZ[263], b11_OFWNT9L_8tZ[262], 
        b11_OFWNT9L_8tZ[261], b11_OFWNT9L_8tZ[260], 
        b11_OFWNT9L_8tZ[259], b11_OFWNT9L_8tZ[258], 
        b11_OFWNT9L_8tZ[257], b11_OFWNT9L_8tZ[256], 
        b11_OFWNT9L_8tZ[255], b11_OFWNT9L_8tZ[254], 
        b11_OFWNT9L_8tZ[253], b11_OFWNT9L_8tZ[252], 
        b11_OFWNT9L_8tZ[251], b11_OFWNT9L_8tZ[250], 
        b11_OFWNT9L_8tZ[249], b11_OFWNT9L_8tZ[248], 
        b11_OFWNT9L_8tZ[247], b11_OFWNT9L_8tZ[246], 
        b11_OFWNT9L_8tZ[245], b11_OFWNT9L_8tZ[244], 
        b11_OFWNT9L_8tZ[243], b11_OFWNT9L_8tZ[242], 
        b11_OFWNT9L_8tZ[241], b11_OFWNT9L_8tZ[240], 
        b11_OFWNT9L_8tZ[239], b11_OFWNT9L_8tZ[238], 
        b11_OFWNT9L_8tZ[237], b11_OFWNT9L_8tZ[236], 
        b11_OFWNT9L_8tZ[235], b11_OFWNT9L_8tZ[234], 
        b11_OFWNT9L_8tZ[233], b11_OFWNT9L_8tZ[232], 
        b11_OFWNT9L_8tZ[231], b11_OFWNT9L_8tZ[230], 
        b11_OFWNT9L_8tZ[229], b11_OFWNT9L_8tZ[228], 
        b11_OFWNT9L_8tZ[227], b11_OFWNT9L_8tZ[226], 
        b11_OFWNT9L_8tZ[225], b11_OFWNT9L_8tZ[224], 
        b11_OFWNT9L_8tZ[223], b11_OFWNT9L_8tZ[222], 
        b11_OFWNT9L_8tZ[221], b11_OFWNT9L_8tZ[220], 
        b11_OFWNT9L_8tZ[219], b11_OFWNT9L_8tZ[218], 
        b11_OFWNT9L_8tZ[217], b11_OFWNT9L_8tZ[216], 
        b11_OFWNT9L_8tZ[215], b11_OFWNT9L_8tZ[214], 
        b11_OFWNT9L_8tZ[213], b11_OFWNT9L_8tZ[212], 
        b11_OFWNT9L_8tZ[211], b11_OFWNT9L_8tZ[210], 
        b11_OFWNT9L_8tZ[209], b11_OFWNT9L_8tZ[208], 
        b11_OFWNT9L_8tZ[207], b11_OFWNT9L_8tZ[206], 
        b11_OFWNT9L_8tZ[205], b11_OFWNT9L_8tZ[204], 
        b11_OFWNT9L_8tZ[203], b11_OFWNT9L_8tZ[202], 
        b11_OFWNT9L_8tZ[201], b11_OFWNT9L_8tZ[200], 
        b11_OFWNT9L_8tZ[199], b11_OFWNT9L_8tZ[198], 
        b11_OFWNT9L_8tZ[197], b11_OFWNT9L_8tZ[196], 
        b11_OFWNT9L_8tZ[195], b11_OFWNT9L_8tZ[194], 
        b11_OFWNT9L_8tZ[193], b11_OFWNT9L_8tZ[192], 
        b11_OFWNT9L_8tZ[191], b11_OFWNT9L_8tZ[190], 
        b11_OFWNT9L_8tZ[189], b11_OFWNT9L_8tZ[188], 
        b11_OFWNT9L_8tZ[187], b11_OFWNT9L_8tZ[186], 
        b11_OFWNT9L_8tZ[185], b11_OFWNT9L_8tZ[184], 
        b11_OFWNT9L_8tZ[183], b11_OFWNT9L_8tZ[182], 
        b11_OFWNT9L_8tZ[181], b11_OFWNT9L_8tZ[180], 
        b11_OFWNT9L_8tZ[179], b11_OFWNT9L_8tZ[178], 
        b11_OFWNT9L_8tZ[177], b11_OFWNT9L_8tZ[176], 
        b11_OFWNT9L_8tZ[175], b11_OFWNT9L_8tZ[174], 
        b11_OFWNT9L_8tZ[173], b11_OFWNT9L_8tZ[172], 
        b11_OFWNT9L_8tZ[171], b11_OFWNT9L_8tZ[170], 
        b11_OFWNT9L_8tZ[169], b11_OFWNT9L_8tZ[168], 
        b11_OFWNT9L_8tZ[167], b11_OFWNT9L_8tZ[166], 
        b11_OFWNT9L_8tZ[165], b11_OFWNT9L_8tZ[164], 
        b11_OFWNT9L_8tZ[163], b11_OFWNT9L_8tZ[162], 
        b11_OFWNT9L_8tZ[161], b11_OFWNT9L_8tZ[160], 
        b11_OFWNT9L_8tZ[159], b11_OFWNT9L_8tZ[158], 
        b11_OFWNT9L_8tZ[157], b11_OFWNT9L_8tZ[156], 
        b11_OFWNT9L_8tZ[155], b11_OFWNT9L_8tZ[154], 
        b11_OFWNT9L_8tZ[153], b11_OFWNT9L_8tZ[152], 
        b11_OFWNT9L_8tZ[151], b11_OFWNT9L_8tZ[150], 
        b11_OFWNT9L_8tZ[149], b11_OFWNT9L_8tZ[148], 
        b11_OFWNT9L_8tZ[147], b11_OFWNT9L_8tZ[146], 
        b11_OFWNT9L_8tZ[145], b11_OFWNT9L_8tZ[144], 
        b11_OFWNT9L_8tZ[143], b11_OFWNT9L_8tZ[142], 
        b11_OFWNT9L_8tZ[141], b11_OFWNT9L_8tZ[140], 
        b11_OFWNT9L_8tZ[139], b11_OFWNT9L_8tZ[138], 
        b11_OFWNT9L_8tZ[137], b11_OFWNT9L_8tZ[136], 
        b11_OFWNT9L_8tZ[135], b11_OFWNT9L_8tZ[134], 
        b11_OFWNT9L_8tZ[133], b11_OFWNT9L_8tZ[132], 
        b11_OFWNT9L_8tZ[131], b11_OFWNT9L_8tZ[130], 
        b11_OFWNT9L_8tZ[129], b11_OFWNT9L_8tZ[128], 
        b11_OFWNT9L_8tZ[127], b11_OFWNT9L_8tZ[126], 
        b11_OFWNT9L_8tZ[125], b11_OFWNT9L_8tZ[124], 
        b11_OFWNT9L_8tZ[123], b11_OFWNT9L_8tZ[122], 
        b11_OFWNT9L_8tZ[121], b11_OFWNT9L_8tZ[120], 
        b11_OFWNT9L_8tZ[119], b11_OFWNT9L_8tZ[118], 
        b11_OFWNT9L_8tZ[117], b11_OFWNT9L_8tZ[116], 
        b11_OFWNT9L_8tZ[115], b11_OFWNT9L_8tZ[114], 
        b11_OFWNT9L_8tZ[113], b11_OFWNT9L_8tZ[112], 
        b11_OFWNT9L_8tZ[111], b11_OFWNT9L_8tZ[110], 
        b11_OFWNT9L_8tZ[109], b11_OFWNT9L_8tZ[108], 
        b11_OFWNT9L_8tZ[107], b11_OFWNT9L_8tZ[106], 
        b11_OFWNT9L_8tZ[105], b11_OFWNT9L_8tZ[104], 
        b11_OFWNT9L_8tZ[103], b11_OFWNT9L_8tZ[102], 
        b11_OFWNT9L_8tZ[101], b11_OFWNT9L_8tZ[100], 
        b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], b11_OFWNT9L_8tZ[97], 
        b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], b11_OFWNT9L_8tZ[94], 
        b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], b11_OFWNT9L_8tZ[91], 
        b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], b11_OFWNT9L_8tZ[88], 
        b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], b11_OFWNT9L_8tZ[85], 
        b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], b11_OFWNT9L_8tZ[82], 
        b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], b11_OFWNT9L_8tZ[79], 
        b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], b11_OFWNT9L_8tZ[76], 
        b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], b11_OFWNT9L_8tZ[73], 
        b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], b11_OFWNT9L_8tZ[70], 
        b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], b11_OFWNT9L_8tZ[67], 
        b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], b11_OFWNT9L_8tZ[64], 
        b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], b11_OFWNT9L_8tZ[61], 
        b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], b11_OFWNT9L_8tZ[58], 
        b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], b11_OFWNT9L_8tZ[55], 
        b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], b11_OFWNT9L_8tZ[52], 
        b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], b11_OFWNT9L_8tZ[49], 
        b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], b11_OFWNT9L_8tZ[46], 
        b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], b11_OFWNT9L_8tZ[43], 
        b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], b11_OFWNT9L_8tZ[40], 
        b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], b11_OFWNT9L_8tZ[37], 
        b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], b11_OFWNT9L_8tZ[34], 
        b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], b11_OFWNT9L_8tZ[31], 
        b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], b11_OFWNT9L_8tZ[28], 
        b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], b11_OFWNT9L_8tZ[25], 
        b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], b11_OFWNT9L_8tZ[22], 
        b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], b11_OFWNT9L_8tZ[19], 
        b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], b11_OFWNT9L_8tZ[16], 
        b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], b11_OFWNT9L_8tZ[13], 
        b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], b11_OFWNT9L_8tZ[10], 
        b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], b11_OFWNT9L_8tZ[7], 
        b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], b11_OFWNT9L_8tZ[4], 
        b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], b11_OFWNT9L_8tZ[1], 
        b11_OFWNT9L_8tZ[0]}), .IICE_comm2iice({IICE_comm2iice[11], 
        IICE_comm2iice[10]}), .b11_PSyil9s_FMZ(b11_PSyil9s_FMZ), 
        .BW_clk_c(BW_clk_c), .b7_PSyi3wy(b7_PSyi3wy), .b4_PLyF(b4_PLyF)
        , .b8_PSyiBgYG(b8_PSyiBgYG));
    GND GND (.Y(GND_net_1));
    b7_OCByLXC_Z1_x_0 b5_nUTGT (.b6_Ocm0rW_0_0_o2({b6_Ocm0rW_0_0_o2[2]})
        , .IICE_comm2iice({IICE_comm2iice[11], IICE_comm2iice[10], 
        IICE_comm2iice[9], IICE_comm2iice[8]}), .b13_nAzGfFM_sLsv3_0(
        b13_nAzGfFM_sLsv3[1]), .b8_SoWGfWYY(b8_SoWGfWYY), 
        .b8_SoWGfWYY_i(b8_SoWGfWYY_i), .BW_clk_c(BW_clk_c), 
        .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh), .b11_PSyil9s_FMZ(
        b11_PSyil9s_FMZ), .b11_uRrc2XfY_XH(b11_uRrc2XfY_XH), .b4_PLyF(
        b4_PLyF), .b13_nUTQBgfDb_Z4D(b13_nUTQBgfDb_Z4D), 
        .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), .b16_nYhI39swMeEd_A78(
        b16_nYhI39swMeEd_A78), .b15_nYhI39swMeEd_Mg(
        b15_nYhI39swMeEd_Mg), .b12_vABZ3qsY_Lyh(b12_vABZ3qsY_Lyh), 
        .b11_vABZ3qsY_XH(b11_vABZ3qsY_XH));
    
endmodule


module b19_nczQ_DYg_YFaRM_oUoP_24s_1s_x_0(
       b12_PSyi_KyDbLbb,
       b8_FZFFLXYE,
       IICE_comm2iice_6,
       IICE_comm2iice_4,
       IICE_comm2iice_5,
       IICE_comm2iice_0,
       IICE_comm2iice_1,
       ttdo,
       un1_b5_OvyH3,
       b8_jAA_KlCO,
       N_21
    );
input  [9:0] b12_PSyi_KyDbLbb;
input  [9:0] b8_FZFFLXYE;
input  IICE_comm2iice_6;
input  IICE_comm2iice_4;
input  IICE_comm2iice_5;
input  IICE_comm2iice_0;
input  IICE_comm2iice_1;
output ttdo;
output un1_b5_OvyH3;
input  b8_jAA_KlCO;
input  N_21;

    wire \b13_PLF_2grFt_FH9[22] , VCC_net_1, 
        \b13_PLF_2grFt_FH9_10[22] , N_14, GND_net_1, 
        \b13_PLF_2grFt_FH9[23] , \b13_PLF_2grFt_FH9_10[23] , 
        \b13_PLF_2grFt_FH9[7] , \b13_PLF_2grFt_FH9_10[7] , 
        \b13_PLF_2grFt_FH9[8] , \b13_PLF_2grFt_FH9_10[8] , 
        \b13_PLF_2grFt_FH9[9] , \b13_PLF_2grFt_FH9_10[9] , 
        \b13_PLF_2grFt_FH9[10] , \b13_PLF_2grFt_FH9_10[10] , 
        \b13_PLF_2grFt_FH9[11] , \b13_PLF_2grFt_FH9_10[11] , 
        \b13_PLF_2grFt_FH9[12] , \b13_PLF_2grFt_FH9_10[12] , 
        \b13_PLF_2grFt_FH9[13] , \b13_PLF_2grFt_FH9_10[13] , 
        \b13_PLF_2grFt_FH9[14] , \b13_PLF_2grFt_FH9_10[14] , 
        \b13_PLF_2grFt_FH9[15] , \b13_PLF_2grFt_FH9_10[15] , 
        \b13_PLF_2grFt_FH9[16] , \b13_PLF_2grFt_FH9_10[16] , 
        \b13_PLF_2grFt_FH9[17] , \b13_PLF_2grFt_FH9_10[17] , 
        \b13_PLF_2grFt_FH9[18] , \b13_PLF_2grFt_FH9_10[18] , 
        \b13_PLF_2grFt_FH9[19] , \b13_PLF_2grFt_FH9_10[19] , 
        \b13_PLF_2grFt_FH9[20] , \b13_PLF_2grFt_FH9_10[20] , 
        \b13_PLF_2grFt_FH9[21] , \b13_PLF_2grFt_FH9_10[21] , 
        \b13_PLF_2grFt_FH9_10[0] , \b13_PLF_2grFt_FH9[1] , 
        \b13_PLF_2grFt_FH9_10[1] , \b13_PLF_2grFt_FH9[2] , 
        \b13_PLF_2grFt_FH9_10[2] , \b13_PLF_2grFt_FH9[3] , 
        \b13_PLF_2grFt_FH9_10[3] , \b13_PLF_2grFt_FH9[4] , 
        \b13_PLF_2grFt_FH9_10[4] , \b13_PLF_2grFt_FH9[5] , 
        \b13_PLF_2grFt_FH9_10[5] , \b13_PLF_2grFt_FH9[6] , 
        \b13_PLF_2grFt_FH9_10[6] ;
    
    CFG2 #( .INIT(4'hE) )  \genblk1.un1_b5_OvyH3  (.A(IICE_comm2iice_4)
        , .B(IICE_comm2iice_5), .Y(un1_b5_OvyH3));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_10[0]  (.A(
        IICE_comm2iice_4), .B(\b13_PLF_2grFt_FH9[1] ), .Y(
        \b13_PLF_2grFt_FH9_10[0] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[19]  (.A(
        b12_PSyi_KyDbLbb[5]), .B(\b13_PLF_2grFt_FH9[20] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[19] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[2]  (.D(\b13_PLF_2grFt_FH9_10[2] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[2] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[22]  (.A(
        b12_PSyi_KyDbLbb[8]), .B(\b13_PLF_2grFt_FH9[23] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[22] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[15]  (.A(
        b12_PSyi_KyDbLbb[1]), .B(\b13_PLF_2grFt_FH9[16] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[15] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[2]  (.A(
        b8_jAA_KlCO), .B(\b13_PLF_2grFt_FH9[3] ), .C(IICE_comm2iice_4), 
        .Y(\b13_PLF_2grFt_FH9_10[2] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[5]  (.D(\b13_PLF_2grFt_FH9_10[5] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[5] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[5]  (.A(
        b8_FZFFLXYE[1]), .B(\b13_PLF_2grFt_FH9[6] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[5] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[16]  (.D(\b13_PLF_2grFt_FH9_10[16] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[16] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_10[1]  (.A(
        IICE_comm2iice_4), .B(\b13_PLF_2grFt_FH9[2] ), .Y(
        \b13_PLF_2grFt_FH9_10[1] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_10[3]  (.A(
        IICE_comm2iice_4), .B(\b13_PLF_2grFt_FH9[4] ), .Y(
        \b13_PLF_2grFt_FH9_10[3] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[10]  (.D(\b13_PLF_2grFt_FH9_10[10] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[10] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[12]  (.A(
        b8_FZFFLXYE[8]), .B(\b13_PLF_2grFt_FH9[13] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[12] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[23]  (.D(\b13_PLF_2grFt_FH9_10[23] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[0]  (.D(\b13_PLF_2grFt_FH9_10[0] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(ttdo));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[6]  (.A(
        b8_FZFFLXYE[2]), .B(\b13_PLF_2grFt_FH9[7] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[6] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[11]  (.D(\b13_PLF_2grFt_FH9_10[11] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[11] ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[9]  (.A(
        b8_FZFFLXYE[5]), .B(\b13_PLF_2grFt_FH9[10] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[12]  (.D(\b13_PLF_2grFt_FH9_10[12] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[12] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[17]  (.D(\b13_PLF_2grFt_FH9_10[17] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[17] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[20]  (.D(\b13_PLF_2grFt_FH9_10[20] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[20] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[14]  (.D(\b13_PLF_2grFt_FH9_10[14] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[14] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[6]  (.D(\b13_PLF_2grFt_FH9_10[6] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[6] ));
    GND GND (.Y(GND_net_1));
    SLE \genblk1.b13_PLF_2grFt_FH9[21]  (.D(\b13_PLF_2grFt_FH9_10[21] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[21] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[17]  (.A(
        b12_PSyi_KyDbLbb[3]), .B(\b13_PLF_2grFt_FH9[18] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[17] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[20]  (.A(
        b12_PSyi_KyDbLbb[6]), .B(\b13_PLF_2grFt_FH9[21] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[20] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[22]  (.D(\b13_PLF_2grFt_FH9_10[22] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[22] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[18]  (.D(\b13_PLF_2grFt_FH9_10[18] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[18] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[21]  (.A(
        b12_PSyi_KyDbLbb[7]), .B(\b13_PLF_2grFt_FH9[22] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[21] ));
    CFG2 #( .INIT(4'h8) )  \genblk1.b13_PLF_2grFt_FH9_10[23]  (.A(
        IICE_comm2iice_4), .B(b12_PSyi_KyDbLbb[9]), .Y(
        \b13_PLF_2grFt_FH9_10[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[9]  (.D(\b13_PLF_2grFt_FH9_10[9] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[4]  (.D(\b13_PLF_2grFt_FH9_10[4] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[4] ));
    CFG4 #( .INIT(16'h8000) )  un1_b13_PLF_2grFt_FH923_i_a2 (.A(
        IICE_comm2iice_0), .B(N_21), .C(IICE_comm2iice_1), .D(
        un1_b5_OvyH3), .Y(N_14));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[10]  (.A(
        b8_FZFFLXYE[6]), .B(\b13_PLF_2grFt_FH9[11] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[10] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[11]  (.A(
        b8_FZFFLXYE[7]), .B(\b13_PLF_2grFt_FH9[12] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[11] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[18]  (.A(
        b12_PSyi_KyDbLbb[4]), .B(\b13_PLF_2grFt_FH9[19] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[18] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[13]  (.A(
        b8_FZFFLXYE[9]), .B(\b13_PLF_2grFt_FH9[14] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[13] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[15]  (.D(\b13_PLF_2grFt_FH9_10[15] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[15] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[3]  (.D(\b13_PLF_2grFt_FH9_10[3] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[3] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[8]  (.A(
        b8_FZFFLXYE[4]), .B(\b13_PLF_2grFt_FH9[9] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[8] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[14]  (.A(
        b12_PSyi_KyDbLbb[0]), .B(\b13_PLF_2grFt_FH9[15] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[14] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[1]  (.D(\b13_PLF_2grFt_FH9_10[1] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[1] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[7]  (.D(\b13_PLF_2grFt_FH9_10[7] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[19]  (.D(\b13_PLF_2grFt_FH9_10[19] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[19] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[7]  (.A(
        b8_FZFFLXYE[3]), .B(\b13_PLF_2grFt_FH9[8] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[8]  (.D(\b13_PLF_2grFt_FH9_10[8] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[8] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[16]  (.A(
        b12_PSyi_KyDbLbb[2]), .B(\b13_PLF_2grFt_FH9[17] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[16] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[4]  (.A(
        b8_FZFFLXYE[0]), .B(\b13_PLF_2grFt_FH9[5] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[4] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[13]  (.D(\b13_PLF_2grFt_FH9_10[13] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[13] ));
    
endmodule


module b13_vFW_xNywD_EdR_383s_10s_1024s_0s_x_0(
       IICE_comm2iice,
       b12_2_St6KCa_jHv,
       b7_vFW_PlM,
       b11_OFWNT9L_8tZ,
       b9_v_mzCDYXs_2,
       b9_v_mzCDYXs_1,
       b9_v_mzCDYXs_0,
       b9_v_mzCDYXs,
       b9_v_mzCDYXs_8,
       b9_v_mzCDYXs_7,
       b9_v_mzCDYXs_6,
       b9_v_mzCDYXs_5,
       b9_v_mzCDYXs_4,
       b9_v_mzCDYXs_3,
       BW_clk_c,
       b4_2o_z
    );
input  [11:11] IICE_comm2iice;
input  [9:0] b12_2_St6KCa_jHv;
output [376:0] b7_vFW_PlM;
input  [376:0] b11_OFWNT9L_8tZ;
input  b9_v_mzCDYXs_2;
input  b9_v_mzCDYXs_1;
input  b9_v_mzCDYXs_0;
input  b9_v_mzCDYXs;
input  b9_v_mzCDYXs_8;
input  b9_v_mzCDYXs_7;
input  b9_v_mzCDYXs_6;
input  b9_v_mzCDYXs_5;
input  b9_v_mzCDYXs_4;
input  b9_v_mzCDYXs_3;
input  BW_clk_c;
input  b4_2o_z;

    wire VCC_net_1, GND_net_1;
    
    RAM1K18 b3_SoW_b3_SoW_0_0 (.A_DOUT({b7_vFW_PlM[17], b7_vFW_PlM[16], 
        b7_vFW_PlM[15], b7_vFW_PlM[14], b7_vFW_PlM[13], b7_vFW_PlM[12], 
        b7_vFW_PlM[11], b7_vFW_PlM[10], b7_vFW_PlM[9], b7_vFW_PlM[8], 
        b7_vFW_PlM[7], b7_vFW_PlM[6], b7_vFW_PlM[5], b7_vFW_PlM[4], 
        b7_vFW_PlM[3], b7_vFW_PlM[2], b7_vFW_PlM[1], b7_vFW_PlM[0]}), 
        .B_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, 
        nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[17], b11_OFWNT9L_8tZ[16], b11_OFWNT9L_8tZ[15], 
        b11_OFWNT9L_8tZ[14], b11_OFWNT9L_8tZ[13], b11_OFWNT9L_8tZ[12], 
        b11_OFWNT9L_8tZ[11], b11_OFWNT9L_8tZ[10], b11_OFWNT9L_8tZ[9], 
        b11_OFWNT9L_8tZ[8], b11_OFWNT9L_8tZ[7], b11_OFWNT9L_8tZ[6], 
        b11_OFWNT9L_8tZ[5], b11_OFWNT9L_8tZ[4], b11_OFWNT9L_8tZ[3], 
        b11_OFWNT9L_8tZ[2], b11_OFWNT9L_8tZ[1], b11_OFWNT9L_8tZ[0]}), 
        .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_6 (.A_DOUT({b7_vFW_PlM[125], 
        b7_vFW_PlM[124], b7_vFW_PlM[123], b7_vFW_PlM[122], 
        b7_vFW_PlM[121], b7_vFW_PlM[120], b7_vFW_PlM[119], 
        b7_vFW_PlM[118], b7_vFW_PlM[117], b7_vFW_PlM[116], 
        b7_vFW_PlM[115], b7_vFW_PlM[114], b7_vFW_PlM[113], 
        b7_vFW_PlM[112], b7_vFW_PlM[111], b7_vFW_PlM[110], 
        b7_vFW_PlM[109], b7_vFW_PlM[108]}), .B_DOUT({nc18, nc19, nc20, 
        nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, nc29, nc30, 
        nc31, nc32, nc33, nc34, nc35}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[125], b11_OFWNT9L_8tZ[124], 
        b11_OFWNT9L_8tZ[123], b11_OFWNT9L_8tZ[122], 
        b11_OFWNT9L_8tZ[121], b11_OFWNT9L_8tZ[120], 
        b11_OFWNT9L_8tZ[119], b11_OFWNT9L_8tZ[118], 
        b11_OFWNT9L_8tZ[117], b11_OFWNT9L_8tZ[116], 
        b11_OFWNT9L_8tZ[115], b11_OFWNT9L_8tZ[114], 
        b11_OFWNT9L_8tZ[113], b11_OFWNT9L_8tZ[112], 
        b11_OFWNT9L_8tZ[111], b11_OFWNT9L_8tZ[110], 
        b11_OFWNT9L_8tZ[109], b11_OFWNT9L_8tZ[108]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_8 (.A_DOUT({b7_vFW_PlM[161], 
        b7_vFW_PlM[160], b7_vFW_PlM[159], b7_vFW_PlM[158], 
        b7_vFW_PlM[157], b7_vFW_PlM[156], b7_vFW_PlM[155], 
        b7_vFW_PlM[154], b7_vFW_PlM[153], b7_vFW_PlM[152], 
        b7_vFW_PlM[151], b7_vFW_PlM[150], b7_vFW_PlM[149], 
        b7_vFW_PlM[148], b7_vFW_PlM[147], b7_vFW_PlM[146], 
        b7_vFW_PlM[145], b7_vFW_PlM[144]}), .B_DOUT({nc36, nc37, nc38, 
        nc39, nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, nc48, 
        nc49, nc50, nc51, nc52, nc53}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[161], b11_OFWNT9L_8tZ[160], 
        b11_OFWNT9L_8tZ[159], b11_OFWNT9L_8tZ[158], 
        b11_OFWNT9L_8tZ[157], b11_OFWNT9L_8tZ[156], 
        b11_OFWNT9L_8tZ[155], b11_OFWNT9L_8tZ[154], 
        b11_OFWNT9L_8tZ[153], b11_OFWNT9L_8tZ[152], 
        b11_OFWNT9L_8tZ[151], b11_OFWNT9L_8tZ[150], 
        b11_OFWNT9L_8tZ[149], b11_OFWNT9L_8tZ[148], 
        b11_OFWNT9L_8tZ[147], b11_OFWNT9L_8tZ[146], 
        b11_OFWNT9L_8tZ[145], b11_OFWNT9L_8tZ[144]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_16 (.A_DOUT({b7_vFW_PlM[305], 
        b7_vFW_PlM[304], b7_vFW_PlM[303], b7_vFW_PlM[302], 
        b7_vFW_PlM[301], b7_vFW_PlM[300], b7_vFW_PlM[299], 
        b7_vFW_PlM[298], b7_vFW_PlM[297], b7_vFW_PlM[296], 
        b7_vFW_PlM[295], b7_vFW_PlM[294], b7_vFW_PlM[293], 
        b7_vFW_PlM[292], b7_vFW_PlM[291], b7_vFW_PlM[290], 
        b7_vFW_PlM[289], b7_vFW_PlM[288]}), .B_DOUT({nc54, nc55, nc56, 
        nc57, nc58, nc59, nc60, nc61, nc62, nc63, nc64, nc65, nc66, 
        nc67, nc68, nc69, nc70, nc71}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[305], b11_OFWNT9L_8tZ[304], 
        b11_OFWNT9L_8tZ[303], b11_OFWNT9L_8tZ[302], 
        b11_OFWNT9L_8tZ[301], b11_OFWNT9L_8tZ[300], 
        b11_OFWNT9L_8tZ[299], b11_OFWNT9L_8tZ[298], 
        b11_OFWNT9L_8tZ[297], b11_OFWNT9L_8tZ[296], 
        b11_OFWNT9L_8tZ[295], b11_OFWNT9L_8tZ[294], 
        b11_OFWNT9L_8tZ[293], b11_OFWNT9L_8tZ[292], 
        b11_OFWNT9L_8tZ[291], b11_OFWNT9L_8tZ[290], 
        b11_OFWNT9L_8tZ[289], b11_OFWNT9L_8tZ[288]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_13 (.A_DOUT({b7_vFW_PlM[251], 
        b7_vFW_PlM[250], b7_vFW_PlM[249], b7_vFW_PlM[248], 
        b7_vFW_PlM[247], b7_vFW_PlM[246], b7_vFW_PlM[245], 
        b7_vFW_PlM[244], b7_vFW_PlM[243], b7_vFW_PlM[242], 
        b7_vFW_PlM[241], b7_vFW_PlM[240], b7_vFW_PlM[239], 
        b7_vFW_PlM[238], b7_vFW_PlM[237], b7_vFW_PlM[236], 
        b7_vFW_PlM[235], b7_vFW_PlM[234]}), .B_DOUT({nc72, nc73, nc74, 
        nc75, nc76, nc77, nc78, nc79, nc80, nc81, nc82, nc83, nc84, 
        nc85, nc86, nc87, nc88, nc89}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[251], b11_OFWNT9L_8tZ[250], 
        b11_OFWNT9L_8tZ[249], b11_OFWNT9L_8tZ[248], 
        b11_OFWNT9L_8tZ[247], b11_OFWNT9L_8tZ[246], 
        b11_OFWNT9L_8tZ[245], b11_OFWNT9L_8tZ[244], 
        b11_OFWNT9L_8tZ[243], b11_OFWNT9L_8tZ[242], 
        b11_OFWNT9L_8tZ[241], b11_OFWNT9L_8tZ[240], 
        b11_OFWNT9L_8tZ[239], b11_OFWNT9L_8tZ[238], 
        b11_OFWNT9L_8tZ[237], b11_OFWNT9L_8tZ[236], 
        b11_OFWNT9L_8tZ[235], b11_OFWNT9L_8tZ[234]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    GND GND (.Y(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_4 (.A_DOUT({b7_vFW_PlM[89], b7_vFW_PlM[88], 
        b7_vFW_PlM[87], b7_vFW_PlM[86], b7_vFW_PlM[85], b7_vFW_PlM[84], 
        b7_vFW_PlM[83], b7_vFW_PlM[82], b7_vFW_PlM[81], b7_vFW_PlM[80], 
        b7_vFW_PlM[79], b7_vFW_PlM[78], b7_vFW_PlM[77], b7_vFW_PlM[76], 
        b7_vFW_PlM[75], b7_vFW_PlM[74], b7_vFW_PlM[73], b7_vFW_PlM[72]})
        , .B_DOUT({nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97, 
        nc98, nc99, nc100, nc101, nc102, nc103, nc104, nc105, nc106, 
        nc107}), .BUSY(), .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(
        IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), 
        .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[89], b11_OFWNT9L_8tZ[88], b11_OFWNT9L_8tZ[87], 
        b11_OFWNT9L_8tZ[86], b11_OFWNT9L_8tZ[85], b11_OFWNT9L_8tZ[84], 
        b11_OFWNT9L_8tZ[83], b11_OFWNT9L_8tZ[82], b11_OFWNT9L_8tZ[81], 
        b11_OFWNT9L_8tZ[80], b11_OFWNT9L_8tZ[79], b11_OFWNT9L_8tZ[78], 
        b11_OFWNT9L_8tZ[77], b11_OFWNT9L_8tZ[76], b11_OFWNT9L_8tZ[75], 
        b11_OFWNT9L_8tZ[74], b11_OFWNT9L_8tZ[73], b11_OFWNT9L_8tZ[72]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_15 (.A_DOUT({b7_vFW_PlM[287], 
        b7_vFW_PlM[286], b7_vFW_PlM[285], b7_vFW_PlM[284], 
        b7_vFW_PlM[283], b7_vFW_PlM[282], b7_vFW_PlM[281], 
        b7_vFW_PlM[280], b7_vFW_PlM[279], b7_vFW_PlM[278], 
        b7_vFW_PlM[277], b7_vFW_PlM[276], b7_vFW_PlM[275], 
        b7_vFW_PlM[274], b7_vFW_PlM[273], b7_vFW_PlM[272], 
        b7_vFW_PlM[271], b7_vFW_PlM[270]}), .B_DOUT({nc108, nc109, 
        nc110, nc111, nc112, nc113, nc114, nc115, nc116, nc117, nc118, 
        nc119, nc120, nc121, nc122, nc123, nc124, nc125}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[287], b11_OFWNT9L_8tZ[286], 
        b11_OFWNT9L_8tZ[285], b11_OFWNT9L_8tZ[284], 
        b11_OFWNT9L_8tZ[283], b11_OFWNT9L_8tZ[282], 
        b11_OFWNT9L_8tZ[281], b11_OFWNT9L_8tZ[280], 
        b11_OFWNT9L_8tZ[279], b11_OFWNT9L_8tZ[278], 
        b11_OFWNT9L_8tZ[277], b11_OFWNT9L_8tZ[276], 
        b11_OFWNT9L_8tZ[275], b11_OFWNT9L_8tZ[274], 
        b11_OFWNT9L_8tZ[273], b11_OFWNT9L_8tZ[272], 
        b11_OFWNT9L_8tZ[271], b11_OFWNT9L_8tZ[270]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_5 (.A_DOUT({b7_vFW_PlM[107], 
        b7_vFW_PlM[106], b7_vFW_PlM[105], b7_vFW_PlM[104], 
        b7_vFW_PlM[103], b7_vFW_PlM[102], b7_vFW_PlM[101], 
        b7_vFW_PlM[100], b7_vFW_PlM[99], b7_vFW_PlM[98], 
        b7_vFW_PlM[97], b7_vFW_PlM[96], b7_vFW_PlM[95], b7_vFW_PlM[94], 
        b7_vFW_PlM[93], b7_vFW_PlM[92], b7_vFW_PlM[91], b7_vFW_PlM[90]})
        , .B_DOUT({nc126, nc127, nc128, nc129, nc130, nc131, nc132, 
        nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, nc141, 
        nc142, nc143}), .BUSY(), .A_CLK(IICE_comm2iice[11]), 
        .A_DOUT_CLK(IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), 
        .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1})
        , .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[107], b11_OFWNT9L_8tZ[106], 
        b11_OFWNT9L_8tZ[105], b11_OFWNT9L_8tZ[104], 
        b11_OFWNT9L_8tZ[103], b11_OFWNT9L_8tZ[102], 
        b11_OFWNT9L_8tZ[101], b11_OFWNT9L_8tZ[100], 
        b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], b11_OFWNT9L_8tZ[97], 
        b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], b11_OFWNT9L_8tZ[94], 
        b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], b11_OFWNT9L_8tZ[91], 
        b11_OFWNT9L_8tZ[90]}), .B_ADDR({b12_2_St6KCa_jHv[9], 
        b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], 
        b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], 
        b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, 
        b4_2o_z}), .A_EN(VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({
        VCC_net_1, GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(
        VCC_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(
        GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_1 (.A_DOUT({b7_vFW_PlM[35], b7_vFW_PlM[34], 
        b7_vFW_PlM[33], b7_vFW_PlM[32], b7_vFW_PlM[31], b7_vFW_PlM[30], 
        b7_vFW_PlM[29], b7_vFW_PlM[28], b7_vFW_PlM[27], b7_vFW_PlM[26], 
        b7_vFW_PlM[25], b7_vFW_PlM[24], b7_vFW_PlM[23], b7_vFW_PlM[22], 
        b7_vFW_PlM[21], b7_vFW_PlM[20], b7_vFW_PlM[19], b7_vFW_PlM[18]})
        , .B_DOUT({nc144, nc145, nc146, nc147, nc148, nc149, nc150, 
        nc151, nc152, nc153, nc154, nc155, nc156, nc157, nc158, nc159, 
        nc160, nc161}), .BUSY(), .A_CLK(IICE_comm2iice[11]), 
        .A_DOUT_CLK(IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), 
        .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1})
        , .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[35], b11_OFWNT9L_8tZ[34], b11_OFWNT9L_8tZ[33], 
        b11_OFWNT9L_8tZ[32], b11_OFWNT9L_8tZ[31], b11_OFWNT9L_8tZ[30], 
        b11_OFWNT9L_8tZ[29], b11_OFWNT9L_8tZ[28], b11_OFWNT9L_8tZ[27], 
        b11_OFWNT9L_8tZ[26], b11_OFWNT9L_8tZ[25], b11_OFWNT9L_8tZ[24], 
        b11_OFWNT9L_8tZ[23], b11_OFWNT9L_8tZ[22], b11_OFWNT9L_8tZ[21], 
        b11_OFWNT9L_8tZ[20], b11_OFWNT9L_8tZ[19], b11_OFWNT9L_8tZ[18]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_3 (.A_DOUT({b7_vFW_PlM[71], b7_vFW_PlM[70], 
        b7_vFW_PlM[69], b7_vFW_PlM[68], b7_vFW_PlM[67], b7_vFW_PlM[66], 
        b7_vFW_PlM[65], b7_vFW_PlM[64], b7_vFW_PlM[63], b7_vFW_PlM[62], 
        b7_vFW_PlM[61], b7_vFW_PlM[60], b7_vFW_PlM[59], b7_vFW_PlM[58], 
        b7_vFW_PlM[57], b7_vFW_PlM[56], b7_vFW_PlM[55], b7_vFW_PlM[54]})
        , .B_DOUT({nc162, nc163, nc164, nc165, nc166, nc167, nc168, 
        nc169, nc170, nc171, nc172, nc173, nc174, nc175, nc176, nc177, 
        nc178, nc179}), .BUSY(), .A_CLK(IICE_comm2iice[11]), 
        .A_DOUT_CLK(IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), 
        .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1})
        , .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[71], b11_OFWNT9L_8tZ[70], b11_OFWNT9L_8tZ[69], 
        b11_OFWNT9L_8tZ[68], b11_OFWNT9L_8tZ[67], b11_OFWNT9L_8tZ[66], 
        b11_OFWNT9L_8tZ[65], b11_OFWNT9L_8tZ[64], b11_OFWNT9L_8tZ[63], 
        b11_OFWNT9L_8tZ[62], b11_OFWNT9L_8tZ[61], b11_OFWNT9L_8tZ[60], 
        b11_OFWNT9L_8tZ[59], b11_OFWNT9L_8tZ[58], b11_OFWNT9L_8tZ[57], 
        b11_OFWNT9L_8tZ[56], b11_OFWNT9L_8tZ[55], b11_OFWNT9L_8tZ[54]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_12 (.A_DOUT({b7_vFW_PlM[233], 
        b7_vFW_PlM[232], b7_vFW_PlM[231], b7_vFW_PlM[230], 
        b7_vFW_PlM[229], b7_vFW_PlM[228], b7_vFW_PlM[227], 
        b7_vFW_PlM[226], b7_vFW_PlM[225], b7_vFW_PlM[224], 
        b7_vFW_PlM[223], b7_vFW_PlM[222], b7_vFW_PlM[221], 
        b7_vFW_PlM[220], b7_vFW_PlM[219], b7_vFW_PlM[218], 
        b7_vFW_PlM[217], b7_vFW_PlM[216]}), .B_DOUT({nc180, nc181, 
        nc182, nc183, nc184, nc185, nc186, nc187, nc188, nc189, nc190, 
        nc191, nc192, nc193, nc194, nc195, nc196, nc197}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[233], b11_OFWNT9L_8tZ[232], 
        b11_OFWNT9L_8tZ[231], b11_OFWNT9L_8tZ[230], 
        b11_OFWNT9L_8tZ[229], b11_OFWNT9L_8tZ[228], 
        b11_OFWNT9L_8tZ[227], b11_OFWNT9L_8tZ[226], 
        b11_OFWNT9L_8tZ[225], b11_OFWNT9L_8tZ[224], 
        b11_OFWNT9L_8tZ[223], b11_OFWNT9L_8tZ[222], 
        b11_OFWNT9L_8tZ[221], b11_OFWNT9L_8tZ[220], 
        b11_OFWNT9L_8tZ[219], b11_OFWNT9L_8tZ[218], 
        b11_OFWNT9L_8tZ[217], b11_OFWNT9L_8tZ[216]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_17 (.A_DOUT({b7_vFW_PlM[323], 
        b7_vFW_PlM[322], b7_vFW_PlM[321], b7_vFW_PlM[320], 
        b7_vFW_PlM[319], b7_vFW_PlM[318], b7_vFW_PlM[317], 
        b7_vFW_PlM[316], b7_vFW_PlM[315], b7_vFW_PlM[314], 
        b7_vFW_PlM[313], b7_vFW_PlM[312], b7_vFW_PlM[311], 
        b7_vFW_PlM[310], b7_vFW_PlM[309], b7_vFW_PlM[308], 
        b7_vFW_PlM[307], b7_vFW_PlM[306]}), .B_DOUT({nc198, nc199, 
        nc200, nc201, nc202, nc203, nc204, nc205, nc206, nc207, nc208, 
        nc209, nc210, nc211, nc212, nc213, nc214, nc215}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[323], b11_OFWNT9L_8tZ[322], 
        b11_OFWNT9L_8tZ[321], b11_OFWNT9L_8tZ[320], 
        b11_OFWNT9L_8tZ[319], b11_OFWNT9L_8tZ[318], 
        b11_OFWNT9L_8tZ[317], b11_OFWNT9L_8tZ[316], 
        b11_OFWNT9L_8tZ[315], b11_OFWNT9L_8tZ[314], 
        b11_OFWNT9L_8tZ[313], b11_OFWNT9L_8tZ[312], 
        b11_OFWNT9L_8tZ[311], b11_OFWNT9L_8tZ[310], 
        b11_OFWNT9L_8tZ[309], b11_OFWNT9L_8tZ[308], 
        b11_OFWNT9L_8tZ[307], b11_OFWNT9L_8tZ[306]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_2 (.A_DOUT({b7_vFW_PlM[53], b7_vFW_PlM[52], 
        b7_vFW_PlM[51], b7_vFW_PlM[50], b7_vFW_PlM[49], b7_vFW_PlM[48], 
        b7_vFW_PlM[47], b7_vFW_PlM[46], b7_vFW_PlM[45], b7_vFW_PlM[44], 
        b7_vFW_PlM[43], b7_vFW_PlM[42], b7_vFW_PlM[41], b7_vFW_PlM[40], 
        b7_vFW_PlM[39], b7_vFW_PlM[38], b7_vFW_PlM[37], b7_vFW_PlM[36]})
        , .B_DOUT({nc216, nc217, nc218, nc219, nc220, nc221, nc222, 
        nc223, nc224, nc225, nc226, nc227, nc228, nc229, nc230, nc231, 
        nc232, nc233}), .BUSY(), .A_CLK(IICE_comm2iice[11]), 
        .A_DOUT_CLK(IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), 
        .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1})
        , .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[53], b11_OFWNT9L_8tZ[52], b11_OFWNT9L_8tZ[51], 
        b11_OFWNT9L_8tZ[50], b11_OFWNT9L_8tZ[49], b11_OFWNT9L_8tZ[48], 
        b11_OFWNT9L_8tZ[47], b11_OFWNT9L_8tZ[46], b11_OFWNT9L_8tZ[45], 
        b11_OFWNT9L_8tZ[44], b11_OFWNT9L_8tZ[43], b11_OFWNT9L_8tZ[42], 
        b11_OFWNT9L_8tZ[41], b11_OFWNT9L_8tZ[40], b11_OFWNT9L_8tZ[39], 
        b11_OFWNT9L_8tZ[38], b11_OFWNT9L_8tZ[37], b11_OFWNT9L_8tZ[36]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_14 (.A_DOUT({b7_vFW_PlM[269], 
        b7_vFW_PlM[268], b7_vFW_PlM[267], b7_vFW_PlM[266], 
        b7_vFW_PlM[265], b7_vFW_PlM[264], b7_vFW_PlM[263], 
        b7_vFW_PlM[262], b7_vFW_PlM[261], b7_vFW_PlM[260], 
        b7_vFW_PlM[259], b7_vFW_PlM[258], b7_vFW_PlM[257], 
        b7_vFW_PlM[256], b7_vFW_PlM[255], b7_vFW_PlM[254], 
        b7_vFW_PlM[253], b7_vFW_PlM[252]}), .B_DOUT({nc234, nc235, 
        nc236, nc237, nc238, nc239, nc240, nc241, nc242, nc243, nc244, 
        nc245, nc246, nc247, nc248, nc249, nc250, nc251}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[269], b11_OFWNT9L_8tZ[268], 
        b11_OFWNT9L_8tZ[267], b11_OFWNT9L_8tZ[266], 
        b11_OFWNT9L_8tZ[265], b11_OFWNT9L_8tZ[264], 
        b11_OFWNT9L_8tZ[263], b11_OFWNT9L_8tZ[262], 
        b11_OFWNT9L_8tZ[261], b11_OFWNT9L_8tZ[260], 
        b11_OFWNT9L_8tZ[259], b11_OFWNT9L_8tZ[258], 
        b11_OFWNT9L_8tZ[257], b11_OFWNT9L_8tZ[256], 
        b11_OFWNT9L_8tZ[255], b11_OFWNT9L_8tZ[254], 
        b11_OFWNT9L_8tZ[253], b11_OFWNT9L_8tZ[252]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_11 (.A_DOUT({b7_vFW_PlM[215], 
        b7_vFW_PlM[214], b7_vFW_PlM[213], b7_vFW_PlM[212], 
        b7_vFW_PlM[211], b7_vFW_PlM[210], b7_vFW_PlM[209], 
        b7_vFW_PlM[208], b7_vFW_PlM[207], b7_vFW_PlM[206], 
        b7_vFW_PlM[205], b7_vFW_PlM[204], b7_vFW_PlM[203], 
        b7_vFW_PlM[202], b7_vFW_PlM[201], b7_vFW_PlM[200], 
        b7_vFW_PlM[199], b7_vFW_PlM[198]}), .B_DOUT({nc252, nc253, 
        nc254, nc255, nc256, nc257, nc258, nc259, nc260, nc261, nc262, 
        nc263, nc264, nc265, nc266, nc267, nc268, nc269}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[215], b11_OFWNT9L_8tZ[214], 
        b11_OFWNT9L_8tZ[213], b11_OFWNT9L_8tZ[212], 
        b11_OFWNT9L_8tZ[211], b11_OFWNT9L_8tZ[210], 
        b11_OFWNT9L_8tZ[209], b11_OFWNT9L_8tZ[208], 
        b11_OFWNT9L_8tZ[207], b11_OFWNT9L_8tZ[206], 
        b11_OFWNT9L_8tZ[205], b11_OFWNT9L_8tZ[204], 
        b11_OFWNT9L_8tZ[203], b11_OFWNT9L_8tZ[202], 
        b11_OFWNT9L_8tZ[201], b11_OFWNT9L_8tZ[200], 
        b11_OFWNT9L_8tZ[199], b11_OFWNT9L_8tZ[198]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_9 (.A_DOUT({b7_vFW_PlM[179], 
        b7_vFW_PlM[178], b7_vFW_PlM[177], b7_vFW_PlM[176], 
        b7_vFW_PlM[175], b7_vFW_PlM[174], b7_vFW_PlM[173], 
        b7_vFW_PlM[172], b7_vFW_PlM[171], b7_vFW_PlM[170], 
        b7_vFW_PlM[169], b7_vFW_PlM[168], b7_vFW_PlM[167], 
        b7_vFW_PlM[166], b7_vFW_PlM[165], b7_vFW_PlM[164], 
        b7_vFW_PlM[163], b7_vFW_PlM[162]}), .B_DOUT({nc270, nc271, 
        nc272, nc273, nc274, nc275, nc276, nc277, nc278, nc279, nc280, 
        nc281, nc282, nc283, nc284, nc285, nc286, nc287}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[179], b11_OFWNT9L_8tZ[178], 
        b11_OFWNT9L_8tZ[177], b11_OFWNT9L_8tZ[176], 
        b11_OFWNT9L_8tZ[175], b11_OFWNT9L_8tZ[174], 
        b11_OFWNT9L_8tZ[173], b11_OFWNT9L_8tZ[172], 
        b11_OFWNT9L_8tZ[171], b11_OFWNT9L_8tZ[170], 
        b11_OFWNT9L_8tZ[169], b11_OFWNT9L_8tZ[168], 
        b11_OFWNT9L_8tZ[167], b11_OFWNT9L_8tZ[166], 
        b11_OFWNT9L_8tZ[165], b11_OFWNT9L_8tZ[164], 
        b11_OFWNT9L_8tZ[163], b11_OFWNT9L_8tZ[162]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_19 (.A_DOUT({b7_vFW_PlM[359], 
        b7_vFW_PlM[358], b7_vFW_PlM[357], b7_vFW_PlM[356], 
        b7_vFW_PlM[355], b7_vFW_PlM[354], b7_vFW_PlM[353], 
        b7_vFW_PlM[352], b7_vFW_PlM[351], b7_vFW_PlM[350], 
        b7_vFW_PlM[349], b7_vFW_PlM[348], b7_vFW_PlM[347], 
        b7_vFW_PlM[346], b7_vFW_PlM[345], b7_vFW_PlM[344], 
        b7_vFW_PlM[343], b7_vFW_PlM[342]}), .B_DOUT({nc288, nc289, 
        nc290, nc291, nc292, nc293, nc294, nc295, nc296, nc297, nc298, 
        nc299, nc300, nc301, nc302, nc303, nc304, nc305}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[359], b11_OFWNT9L_8tZ[358], 
        b11_OFWNT9L_8tZ[357], b11_OFWNT9L_8tZ[356], 
        b11_OFWNT9L_8tZ[355], b11_OFWNT9L_8tZ[354], 
        b11_OFWNT9L_8tZ[353], b11_OFWNT9L_8tZ[352], 
        b11_OFWNT9L_8tZ[351], b11_OFWNT9L_8tZ[350], 
        b11_OFWNT9L_8tZ[349], b11_OFWNT9L_8tZ[348], 
        b11_OFWNT9L_8tZ[347], b11_OFWNT9L_8tZ[346], 
        b11_OFWNT9L_8tZ[345], b11_OFWNT9L_8tZ[344], 
        b11_OFWNT9L_8tZ[343], b11_OFWNT9L_8tZ[342]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_18 (.A_DOUT({b7_vFW_PlM[341], 
        b7_vFW_PlM[340], b7_vFW_PlM[339], b7_vFW_PlM[338], 
        b7_vFW_PlM[337], b7_vFW_PlM[336], b7_vFW_PlM[335], 
        b7_vFW_PlM[334], b7_vFW_PlM[333], b7_vFW_PlM[332], 
        b7_vFW_PlM[331], b7_vFW_PlM[330], b7_vFW_PlM[329], 
        b7_vFW_PlM[328], b7_vFW_PlM[327], b7_vFW_PlM[326], 
        b7_vFW_PlM[325], b7_vFW_PlM[324]}), .B_DOUT({nc306, nc307, 
        nc308, nc309, nc310, nc311, nc312, nc313, nc314, nc315, nc316, 
        nc317, nc318, nc319, nc320, nc321, nc322, nc323}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[341], b11_OFWNT9L_8tZ[340], 
        b11_OFWNT9L_8tZ[339], b11_OFWNT9L_8tZ[338], 
        b11_OFWNT9L_8tZ[337], b11_OFWNT9L_8tZ[336], 
        b11_OFWNT9L_8tZ[335], b11_OFWNT9L_8tZ[334], 
        b11_OFWNT9L_8tZ[333], b11_OFWNT9L_8tZ[332], 
        b11_OFWNT9L_8tZ[331], b11_OFWNT9L_8tZ[330], 
        b11_OFWNT9L_8tZ[329], b11_OFWNT9L_8tZ[328], 
        b11_OFWNT9L_8tZ[327], b11_OFWNT9L_8tZ[326], 
        b11_OFWNT9L_8tZ[325], b11_OFWNT9L_8tZ[324]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_10 (.A_DOUT({b7_vFW_PlM[197], 
        b7_vFW_PlM[196], b7_vFW_PlM[195], b7_vFW_PlM[194], 
        b7_vFW_PlM[193], b7_vFW_PlM[192], b7_vFW_PlM[191], 
        b7_vFW_PlM[190], b7_vFW_PlM[189], b7_vFW_PlM[188], 
        b7_vFW_PlM[187], b7_vFW_PlM[186], b7_vFW_PlM[185], 
        b7_vFW_PlM[184], b7_vFW_PlM[183], b7_vFW_PlM[182], 
        b7_vFW_PlM[181], b7_vFW_PlM[180]}), .B_DOUT({nc324, nc325, 
        nc326, nc327, nc328, nc329, nc330, nc331, nc332, nc333, nc334, 
        nc335, nc336, nc337, nc338, nc339, nc340, nc341}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[197], b11_OFWNT9L_8tZ[196], 
        b11_OFWNT9L_8tZ[195], b11_OFWNT9L_8tZ[194], 
        b11_OFWNT9L_8tZ[193], b11_OFWNT9L_8tZ[192], 
        b11_OFWNT9L_8tZ[191], b11_OFWNT9L_8tZ[190], 
        b11_OFWNT9L_8tZ[189], b11_OFWNT9L_8tZ[188], 
        b11_OFWNT9L_8tZ[187], b11_OFWNT9L_8tZ[186], 
        b11_OFWNT9L_8tZ[185], b11_OFWNT9L_8tZ[184], 
        b11_OFWNT9L_8tZ[183], b11_OFWNT9L_8tZ[182], 
        b11_OFWNT9L_8tZ[181], b11_OFWNT9L_8tZ[180]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_7 (.A_DOUT({b7_vFW_PlM[143], 
        b7_vFW_PlM[142], b7_vFW_PlM[141], b7_vFW_PlM[140], 
        b7_vFW_PlM[139], b7_vFW_PlM[138], b7_vFW_PlM[137], 
        b7_vFW_PlM[136], b7_vFW_PlM[135], b7_vFW_PlM[134], 
        b7_vFW_PlM[133], b7_vFW_PlM[132], b7_vFW_PlM[131], 
        b7_vFW_PlM[130], b7_vFW_PlM[129], b7_vFW_PlM[128], 
        b7_vFW_PlM[127], b7_vFW_PlM[126]}), .B_DOUT({nc342, nc343, 
        nc344, nc345, nc346, nc347, nc348, nc349, nc350, nc351, nc352, 
        nc353, nc354, nc355, nc356, nc357, nc358, nc359}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[143], b11_OFWNT9L_8tZ[142], 
        b11_OFWNT9L_8tZ[141], b11_OFWNT9L_8tZ[140], 
        b11_OFWNT9L_8tZ[139], b11_OFWNT9L_8tZ[138], 
        b11_OFWNT9L_8tZ[137], b11_OFWNT9L_8tZ[136], 
        b11_OFWNT9L_8tZ[135], b11_OFWNT9L_8tZ[134], 
        b11_OFWNT9L_8tZ[133], b11_OFWNT9L_8tZ[132], 
        b11_OFWNT9L_8tZ[131], b11_OFWNT9L_8tZ[130], 
        b11_OFWNT9L_8tZ[129], b11_OFWNT9L_8tZ[128], 
        b11_OFWNT9L_8tZ[127], b11_OFWNT9L_8tZ[126]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_20 (.A_DOUT({nc360, b7_vFW_PlM[376], 
        b7_vFW_PlM[375], b7_vFW_PlM[374], b7_vFW_PlM[373], 
        b7_vFW_PlM[372], b7_vFW_PlM[371], b7_vFW_PlM[370], 
        b7_vFW_PlM[369], b7_vFW_PlM[368], b7_vFW_PlM[367], 
        b7_vFW_PlM[366], b7_vFW_PlM[365], b7_vFW_PlM[364], 
        b7_vFW_PlM[363], b7_vFW_PlM[362], b7_vFW_PlM[361], 
        b7_vFW_PlM[360]}), .B_DOUT({nc361, nc362, nc363, nc364, nc365, 
        nc366, nc367, nc368, nc369, nc370, nc371, nc372, nc373, nc374, 
        nc375, nc376, nc377, nc378}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({GND_net_1, 
        b11_OFWNT9L_8tZ[376], b11_OFWNT9L_8tZ[375], 
        b11_OFWNT9L_8tZ[374], b11_OFWNT9L_8tZ[373], 
        b11_OFWNT9L_8tZ[372], b11_OFWNT9L_8tZ[371], 
        b11_OFWNT9L_8tZ[370], b11_OFWNT9L_8tZ[369], 
        b11_OFWNT9L_8tZ[368], b11_OFWNT9L_8tZ[367], 
        b11_OFWNT9L_8tZ[366], b11_OFWNT9L_8tZ[365], 
        b11_OFWNT9L_8tZ[364], b11_OFWNT9L_8tZ[363], 
        b11_OFWNT9L_8tZ[362], b11_OFWNT9L_8tZ[361], 
        b11_OFWNT9L_8tZ[360]}), .B_ADDR({b12_2_St6KCa_jHv[9], 
        b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], 
        b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], 
        b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, 
        b4_2o_z}), .A_EN(VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({
        VCC_net_1, GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(
        VCC_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(
        GND_net_1));
    
endmodule


module b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0(
       IICE_comm2iice_11,
       IICE_comm2iice_9,
       IICE_comm2iice_1,
       IICE_comm2iice_3,
       IICE_comm2iice_2,
       IICE_comm2iice_4,
       IICE_comm2iice_0,
       IICE_comm2iice_5,
       IICE_comm2iice_6,
       b4_ycsM,
       un1_b13_PLF_2grFt_FH911_i_a2_0_2,
       N_21,
       un1_b5_OvyH3
    );
input  IICE_comm2iice_11;
input  IICE_comm2iice_9;
input  IICE_comm2iice_1;
input  IICE_comm2iice_3;
input  IICE_comm2iice_2;
input  IICE_comm2iice_4;
input  IICE_comm2iice_0;
input  IICE_comm2iice_5;
input  IICE_comm2iice_6;
output b4_ycsM;
output un1_b13_PLF_2grFt_FH911_i_a2_0_2;
output N_21;
input  un1_b5_OvyH3;

    wire \b13_PLF_2grFt_FH9[24] , VCC_net_1, \b13_PLF_2grFt_FH9_5[24] , 
        N_13, GND_net_1, \b13_PLF_2grFt_FH9[25] , 
        \b13_PLF_2grFt_FH9_5[25] , \b13_PLF_2grFt_FH9[26] , 
        \b13_PLF_2grFt_FH9_5[26] , \b13_PLF_2grFt_FH9[27] , 
        \b13_PLF_2grFt_FH9_5[27] , \b13_PLF_2grFt_FH9[28] , 
        \b13_PLF_2grFt_FH9_5[28] , \b13_PLF_2grFt_FH9[29] , 
        \b13_PLF_2grFt_FH9_5[29] , \b13_PLF_2grFt_FH9[30] , 
        \b13_PLF_2grFt_FH9_5[30] , \b13_PLF_2grFt_FH9[31] , 
        \b13_PLF_2grFt_FH9[9] , \b13_PLF_2grFt_FH9_5[9] , 
        \b13_PLF_2grFt_FH9[10] , \b13_PLF_2grFt_FH9_5[10] , 
        \b13_PLF_2grFt_FH9[11] , \b13_PLF_2grFt_FH9_5[11] , 
        \b13_PLF_2grFt_FH9[12] , \b13_PLF_2grFt_FH9_5[12] , 
        \b13_PLF_2grFt_FH9[13] , \b13_PLF_2grFt_FH9_5[13] , 
        \b13_PLF_2grFt_FH9[14] , \b13_PLF_2grFt_FH9_5[14] , 
        \b13_PLF_2grFt_FH9[15] , \b13_PLF_2grFt_FH9_5[15] , 
        \b13_PLF_2grFt_FH9[16] , \b13_PLF_2grFt_FH9_5[16] , 
        \b13_PLF_2grFt_FH9[17] , \b13_PLF_2grFt_FH9_5[17] , 
        \b13_PLF_2grFt_FH9[18] , \b13_PLF_2grFt_FH9_5[18] , 
        \b13_PLF_2grFt_FH9[19] , \b13_PLF_2grFt_FH9_5[19] , 
        \b13_PLF_2grFt_FH9[20] , \b13_PLF_2grFt_FH9_5[20] , 
        \b13_PLF_2grFt_FH9[21] , \b13_PLF_2grFt_FH9_5[21] , 
        \b13_PLF_2grFt_FH9[22] , \b13_PLF_2grFt_FH9_5[22] , 
        \b13_PLF_2grFt_FH9[23] , \b13_PLF_2grFt_FH9_5[23] , 
        \b13_PLF_2grFt_FH9_5[0] , \b13_PLF_2grFt_FH9[1] , 
        \b13_PLF_2grFt_FH9_5[1] , \b13_PLF_2grFt_FH9[2] , 
        \b13_PLF_2grFt_FH9_5[2] , \b13_PLF_2grFt_FH9[3] , 
        \b13_PLF_2grFt_FH9_5[3] , \b13_PLF_2grFt_FH9[4] , 
        \b13_PLF_2grFt_FH9_5[4] , \b13_PLF_2grFt_FH9[5] , 
        \b13_PLF_2grFt_FH9_5[5] , \b13_PLF_2grFt_FH9[6] , 
        \b13_PLF_2grFt_FH9_5[6] , \b13_PLF_2grFt_FH9[7] , 
        \b13_PLF_2grFt_FH9_5[7] , \b13_PLF_2grFt_FH9[8] , 
        \b13_PLF_2grFt_FH9_5[8] ;
    
    SLE \genblk1.b13_PLF_2grFt_FH9[2]  (.D(\b13_PLF_2grFt_FH9_5[2] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[2] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[22]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[23] ), .Y(
        \b13_PLF_2grFt_FH9_5[22] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[26]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[27] ), .Y(
        \b13_PLF_2grFt_FH9_5[26] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[5]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[6] ), .Y(
        \b13_PLF_2grFt_FH9_5[5] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[5]  (.D(\b13_PLF_2grFt_FH9_5[5] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[5] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[16]  (.D(\b13_PLF_2grFt_FH9_5[16] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[16] ));
    CFG3 #( .INIT(8'h20) )  un1_b13_PLF_2grFt_FH911_i_a2_0_2_inst_1 (
        .A(IICE_comm2iice_1), .B(IICE_comm2iice_3), .C(
        IICE_comm2iice_2), .Y(un1_b13_PLF_2grFt_FH911_i_a2_0_2));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[3]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[4] ), .Y(
        \b13_PLF_2grFt_FH9_5[3] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[10]  (.D(\b13_PLF_2grFt_FH9_5[10] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[10] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[25]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[26] ), .Y(
        \b13_PLF_2grFt_FH9_5[25] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[23]  (.D(\b13_PLF_2grFt_FH9_5[23] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[0]  (.D(\b13_PLF_2grFt_FH9_5[0] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b4_ycsM));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[30]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[31] ), .Y(
        \b13_PLF_2grFt_FH9_5[30] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[20]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[21] ), .Y(
        \b13_PLF_2grFt_FH9_5[20] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[11]  (.D(\b13_PLF_2grFt_FH9_5[11] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[11] ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[21]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[22] ), .Y(
        \b13_PLF_2grFt_FH9_5[21] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[18]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[19] ), .Y(
        \b13_PLF_2grFt_FH9_5[18] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[1]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[2] ), .Y(
        \b13_PLF_2grFt_FH9_5[1] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[12]  (.D(\b13_PLF_2grFt_FH9_5[12] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[12] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[17]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[18] ), .Y(
        \b13_PLF_2grFt_FH9_5[17] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[4]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[5] ), .Y(
        \b13_PLF_2grFt_FH9_5[4] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[17]  (.D(\b13_PLF_2grFt_FH9_5[17] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[17] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[26]  (.D(\b13_PLF_2grFt_FH9_5[26] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[26] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[20]  (.D(\b13_PLF_2grFt_FH9_5[20] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[20] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[24]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[25] ), .Y(
        \b13_PLF_2grFt_FH9_5[24] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[13]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[14] ), .Y(
        \b13_PLF_2grFt_FH9_5[13] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[14]  (.D(\b13_PLF_2grFt_FH9_5[14] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[14] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[29]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[30] ), .Y(
        \b13_PLF_2grFt_FH9_5[29] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[6]  (.D(\b13_PLF_2grFt_FH9_5[6] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[6] ));
    GND GND (.Y(GND_net_1));
    SLE \genblk1.b13_PLF_2grFt_FH9[21]  (.D(\b13_PLF_2grFt_FH9_5[21] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[21] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[0]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[1] ), .Y(
        \b13_PLF_2grFt_FH9_5[0] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[22]  (.D(\b13_PLF_2grFt_FH9_5[22] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[22] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[18]  (.D(\b13_PLF_2grFt_FH9_5[18] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[18] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[12]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[13] ), .Y(
        \b13_PLF_2grFt_FH9_5[12] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[16]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[17] ), .Y(
        \b13_PLF_2grFt_FH9_5[16] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[9]  (.D(\b13_PLF_2grFt_FH9_5[9] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[4]  (.D(\b13_PLF_2grFt_FH9_5[4] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[4] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[27]  (.D(\b13_PLF_2grFt_FH9_5[27] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[27] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[30]  (.D(\b13_PLF_2grFt_FH9_5[30] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[30] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[8]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[9] ), .Y(
        \b13_PLF_2grFt_FH9_5[8] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[24]  (.D(\b13_PLF_2grFt_FH9_5[24] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[24] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[15]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[16] ), .Y(
        \b13_PLF_2grFt_FH9_5[15] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[15]  (.D(\b13_PLF_2grFt_FH9_5[15] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[15] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[10]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[11] ), .Y(
        \b13_PLF_2grFt_FH9_5[10] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[3]  (.D(\b13_PLF_2grFt_FH9_5[3] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[3] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[31]  (.D(IICE_comm2iice_9), .CLK(
        IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_PLF_2grFt_FH9[31] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[9]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[10] ), .Y(
        \b13_PLF_2grFt_FH9_5[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[1]  (.D(\b13_PLF_2grFt_FH9_5[1] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[1] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[11]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[12] ), .Y(
        \b13_PLF_2grFt_FH9_5[11] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[7]  (.D(\b13_PLF_2grFt_FH9_5[7] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[19]  (.D(\b13_PLF_2grFt_FH9_5[19] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[19] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[6]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[7] ), .Y(
        \b13_PLF_2grFt_FH9_5[6] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[7]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[8] ), .Y(
        \b13_PLF_2grFt_FH9_5[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[28]  (.D(\b13_PLF_2grFt_FH9_5[28] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[28] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[28]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[29] ), .Y(
        \b13_PLF_2grFt_FH9_5[28] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[8]  (.D(\b13_PLF_2grFt_FH9_5[8] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[8] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[27]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[28] ), .Y(
        \b13_PLF_2grFt_FH9_5[27] ));
    CFG4 #( .INIT(16'h4000) )  un1_b13_PLF_2grFt_FH911_i_a2 (.A(
        IICE_comm2iice_5), .B(N_21), .C(IICE_comm2iice_6), .D(
        un1_b5_OvyH3), .Y(N_13));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[14]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[15] ), .Y(
        \b13_PLF_2grFt_FH9_5[14] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[2]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[3] ), .Y(
        \b13_PLF_2grFt_FH9_5[2] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[25]  (.D(\b13_PLF_2grFt_FH9_5[25] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[25] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[19]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[20] ), .Y(
        \b13_PLF_2grFt_FH9_5[19] ));
    CFG3 #( .INIT(8'h40) )  un1_b13_PLF_2grFt_FH911_i_a2_0 (.A(
        IICE_comm2iice_4), .B(un1_b13_PLF_2grFt_FH911_i_a2_0_2), .C(
        IICE_comm2iice_0), .Y(N_21));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[23]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[24] ), .Y(
        \b13_PLF_2grFt_FH9_5[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[29]  (.D(\b13_PLF_2grFt_FH9_5[29] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[29] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[13]  (.D(\b13_PLF_2grFt_FH9_5[13] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[13] ));
    
endmodule


module b11_SoWyP0zEFKY_383s_0s_6s_0s_2s_2s_0s_0s_2s_0s_x_0(
       b11_OFWNT9L_8tZ,
       mdiclink_reg,
       b6_Ocm0rW_0_0_o2,
       b13_nAzGfFM_sLsv3,
       BW_clk_c,
       b4_2o_z,
       b8_SoWGfWYY,
       b13_oRB_MqCD2_EdR_RNI9OIA
    );
output [376:0] b11_OFWNT9L_8tZ;
input  [376:0] mdiclink_reg;
input  [2:2] b6_Ocm0rW_0_0_o2;
input  [1:1] b13_nAzGfFM_sLsv3;
input  BW_clk_c;
output b4_2o_z;
input  b8_SoWGfWYY;
output b13_oRB_MqCD2_EdR_RNI9OIA;

    wire VCC_net_1, GND_net_1, b13_oRB_MqCD2_EdR;
    
    SLE \genblk2.b5_oRB_C[337]  (.D(mdiclink_reg[39]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[337]));
    SLE \genblk2.b5_oRB_C[207]  (.D(mdiclink_reg[169]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[207]));
    SLE \genblk2.b5_oRB_C[276]  (.D(mdiclink_reg[100]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[276]));
    SLE \genblk2.b5_oRB_C[338]  (.D(mdiclink_reg[38]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[338]));
    SLE \genblk2.b5_oRB_C[324]  (.D(mdiclink_reg[52]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[324]));
    SLE \genblk2.b5_oRB_C[236]  (.D(mdiclink_reg[140]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[236]));
    SLE \genblk2.b5_oRB_C[72]  (.D(mdiclink_reg[304]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[72]));
    SLE \genblk2.b5_oRB_C[171]  (.D(mdiclink_reg[205]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[171]));
    SLE \genblk2.b5_oRB_C[164]  (.D(mdiclink_reg[212]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[164]));
    SLE \genblk2.b5_oRB_C[61]  (.D(mdiclink_reg[315]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[61]));
    SLE \genblk2.b5_oRB_C[131]  (.D(mdiclink_reg[245]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[131]));
    SLE \genblk2.b5_oRB_C[82]  (.D(mdiclink_reg[294]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[82]));
    SLE \genblk2.b5_oRB_C[122]  (.D(mdiclink_reg[254]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[122]));
    SLE \genblk2.b5_oRB_C[341]  (.D(mdiclink_reg[35]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[341]));
    SLE \genblk2.b5_oRB_C[17]  (.D(mdiclink_reg[359]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[17]));
    SLE \genblk2.b5_oRB_C[219]  (.D(mdiclink_reg[157]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[219]));
    SLE \genblk2.b5_oRB_C[327]  (.D(mdiclink_reg[49]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[327]));
    SLE \genblk2.b5_oRB_C[18]  (.D(mdiclink_reg[358]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[18]));
    SLE \genblk2.b5_oRB_C[241]  (.D(mdiclink_reg[135]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[241]));
    SLE \genblk2.b5_oRB_C[66]  (.D(mdiclink_reg[310]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[66]));
    SLE \genblk2.b5_oRB_C[298]  (.D(mdiclink_reg[78]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[298]));
    SLE \genblk2.b5_oRB_C[177]  (.D(mdiclink_reg[199]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[177]));
    SLE \genblk2.b5_oRB_C[328]  (.D(mdiclink_reg[48]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[328]));
    SLE \genblk2.b5_oRB_C[137]  (.D(mdiclink_reg[239]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[137]));
    SLE \genblk2.b5_oRB_C[226]  (.D(mdiclink_reg[150]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[226]));
    SLE \genblk2.b5_oRB_C[259]  (.D(mdiclink_reg[117]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[259]));
    SLE \genblk2.b5_oRB_C[105]  (.D(mdiclink_reg[271]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[105]));
    SLE \genblk2.b5_oRB_C[121]  (.D(mdiclink_reg[255]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[121]));
    SLE \genblk2.b5_oRB_C[306]  (.D(mdiclink_reg[70]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[306]));
    SLE \genblk2.b5_oRB_C[166]  (.D(mdiclink_reg[210]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[166]));
    SLE \genblk2.b5_oRB_C[20]  (.D(mdiclink_reg[356]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[20]));
    SLE \genblk2.b5_oRB_C[43]  (.D(mdiclink_reg[333]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[43]));
    SLE \genblk2.b5_oRB_C[93]  (.D(mdiclink_reg[283]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[93]));
    SLE \genblk2.b5_oRB_C[313]  (.D(mdiclink_reg[63]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[313]));
    SLE \genblk2.b5_oRB_C[205]  (.D(mdiclink_reg[171]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[205]));
    SLE \genblk2.b5_oRB_C[11]  (.D(mdiclink_reg[365]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[11]));
    SLE \genblk2.b5_oRB_C[127]  (.D(mdiclink_reg[249]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[127]));
    SLE \genblk2.b5_oRB_C[30]  (.D(mdiclink_reg[346]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[30]));
    SLE \genblk2.b5_oRB_C[353]  (.D(mdiclink_reg[23]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[353]));
    SLE \genblk2.b5_oRB_C[370]  (.D(mdiclink_reg[6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[370]));
    SLE \genblk2.b5_oRB_C[203]  (.D(mdiclink_reg[173]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[203]));
    SLE \genblk2.b5_oRB_C[330]  (.D(mdiclink_reg[46]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[330]));
    SLE \genblk2.b5_oRB_C[16]  (.D(mdiclink_reg[360]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[16]));
    SLE \genblk2.b5_oRB_C[45]  (.D(mdiclink_reg[331]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[45]));
    SLE \genblk2.b5_oRB_C[299]  (.D(mdiclink_reg[77]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[299]));
    SLE \genblk2.b5_oRB_C[95]  (.D(mdiclink_reg[281]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[95]));
    SLE \genblk2.b5_oRB_C[287]  (.D(mdiclink_reg[89]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[287]));
    SLE \genblk2.b5_oRB_C[248]  (.D(mdiclink_reg[128]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[248]));
    SLE \genblk2.b5_oRB_C[70]  (.D(mdiclink_reg[306]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[70]));
    SLE \genblk2.b5_oRB_C[5]  (.D(mdiclink_reg[371]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[5]));
    SLE \genblk2.b5_oRB_C[80]  (.D(mdiclink_reg[296]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[80]));
    SLE \genblk2.b5_oRB_C[0]  (.D(mdiclink_reg[376]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[0]));
    SLE \genblk2.b5_oRB_C[104]  (.D(mdiclink_reg[272]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[104]));
    SLE \genblk2.b5_oRB_C[57]  (.D(mdiclink_reg[319]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[57]));
    SLE \genblk2.b5_oRB_C[320]  (.D(mdiclink_reg[56]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[320]));
    SLE \genblk2.b5_oRB_C[58]  (.D(mdiclink_reg[318]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[58]));
    SLE \genblk2.b5_oRB_C[63]  (.D(mdiclink_reg[313]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[63]));
    SLE \genblk2.b5_oRB_C[217]  (.D(mdiclink_reg[159]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[217]));
    SLE \genblk2.b5_oRB_C[260]  (.D(mdiclink_reg[116]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[260]));
    SLE \genblk2.b5_oRB_C[185]  (.D(mdiclink_reg[191]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[185]));
    SLE \genblk2.b5_oRB_C[257]  (.D(mdiclink_reg[119]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[257]));
    SLE \genblk2.b5_oRB_C[264]  (.D(mdiclink_reg[112]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[264]));
    SLE \genblk2.b5_oRB_C[249]  (.D(mdiclink_reg[127]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[249]));
    SLE \genblk2.b5_oRB_C[168]  (.D(mdiclink_reg[208]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[168]));
    SLE \genblk2.b5_oRB_C[106]  (.D(mdiclink_reg[270]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[106]));
    SLE \genblk2.b5_oRB_C[65]  (.D(mdiclink_reg[311]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[65]));
    SLE \genblk2.b5_oRB_C[285]  (.D(mdiclink_reg[91]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[285]));
    GND GND (.Y(GND_net_1));
    SLE \genblk2.b5_oRB_C[51]  (.D(mdiclink_reg[325]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[51]));
    SLE \genblk2.b5_oRB_C[365]  (.D(mdiclink_reg[11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[365]));
    SLE \genblk2.b5_oRB_C[371]  (.D(mdiclink_reg[5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[371]));
    SLE \genblk2.b5_oRB_C[362]  (.D(mdiclink_reg[14]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[362]));
    SLE \genblk2.b5_oRB_C[331]  (.D(mdiclink_reg[45]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[331]));
    SLE \genblk2.b5_oRB_C[115]  (.D(mdiclink_reg[261]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[115]));
    SLE \genblk2.b5_oRB_C[283]  (.D(mdiclink_reg[93]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[283]));
    SLE \genblk2.b5_oRB_C[271]  (.D(mdiclink_reg[105]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[271]));
    SLE \genblk2.b5_oRB_C[13]  (.D(mdiclink_reg[363]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[13]));
    SLE \genblk2.b5_oRB_C[56]  (.D(mdiclink_reg[320]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[56]));
    SLE \genblk2.b5_oRB_C[316]  (.D(mdiclink_reg[60]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[316]));
    SLE \genblk2.b5_oRB_C[231]  (.D(mdiclink_reg[145]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[231]));
    SLE \genblk2.b5_oRB_C[343]  (.D(mdiclink_reg[33]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[343]));
    SLE \genblk2.b5_oRB_C[297]  (.D(mdiclink_reg[79]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[297]));
    SLE \genblk2.b5_oRB_C[262]  (.D(mdiclink_reg[114]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[262]));
    SLE \genblk2.b5_oRB_C[215]  (.D(mdiclink_reg[161]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[215]));
    SLE \genblk2.b5_oRB_C[160]  (.D(mdiclink_reg[216]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[160]));
    SLE \genblk2.b5_oRB_C[155]  (.D(mdiclink_reg[221]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[155]));
    SLE \genblk2.b5_oRB_C[163]  (.D(mdiclink_reg[213]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[163]));
    SLE \genblk2.b5_oRB_C[356]  (.D(mdiclink_reg[20]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[356]));
    SLE \genblk2.b5_oRB_C[44]  (.D(mdiclink_reg[332]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[44]));
    SLE \genblk2.b5_oRB_C[321]  (.D(mdiclink_reg[55]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[321]));
    SLE \genblk2.b5_oRB_C[94]  (.D(mdiclink_reg[282]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[94]));
    SLE \genblk2.b5_oRB_C[255]  (.D(mdiclink_reg[121]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[255]));
    SLE \genblk2.b5_oRB_C[184]  (.D(mdiclink_reg[192]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[184]));
    SLE \genblk2.b5_oRB_C[15]  (.D(mdiclink_reg[361]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[15]));
    SLE \genblk2.b5_oRB_C[221]  (.D(mdiclink_reg[155]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[221]));
    SLE \genblk2.b5_oRB_C[213]  (.D(mdiclink_reg[163]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[213]));
    CFG2 #( .INIT(4'hE) )  \genblk2.b13_oRB_MqCD2_EdR_RNI9OIA  (.A(
        b4_2o_z), .B(b8_SoWGfWYY), .Y(b13_oRB_MqCD2_EdR_RNI9OIA));
    SLE \genblk2.b5_oRB_C[369]  (.D(mdiclink_reg[7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[369]));
    SLE \genblk2.b5_oRB_C[253]  (.D(mdiclink_reg[123]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[253]));
    SLE \genblk2.b5_oRB_C[200]  (.D(mdiclink_reg[176]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[200]));
    SLE \genblk2.b5_oRB_C[3]  (.D(mdiclink_reg[373]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[3]));
    SLE \genblk2.b5_oRB_C[195]  (.D(mdiclink_reg[181]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[195]));
    SLE \genblk2.b5_oRB_C[278]  (.D(mdiclink_reg[98]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[278]));
    SLE \genblk2.b5_oRB_C[186]  (.D(mdiclink_reg[190]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[186]));
    SLE \genblk2.b5_oRB_C[114]  (.D(mdiclink_reg[262]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[114]));
    SLE \genblk2.b5_oRB_C[238]  (.D(mdiclink_reg[138]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[238]));
    SLE \genblk2.b5_oRB_C[204]  (.D(mdiclink_reg[172]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[204]));
    SLE \genblk2.b5_oRB_C[247]  (.D(mdiclink_reg[129]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[247]));
    SLE \genblk2.b5_oRB_C[108]  (.D(mdiclink_reg[268]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[108]));
    SLE \genblk2.b5_oRB_C[295]  (.D(mdiclink_reg[81]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[295]));
    SLE \genblk2.b5_oRB_C[169]  (.D(mdiclink_reg[207]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[169]));
    SLE \genblk2.b5_oRB_C[154]  (.D(mdiclink_reg[222]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[154]));
    SLE \genblk2.b5_oRB_C[305]  (.D(mdiclink_reg[71]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[305]));
    SLE \genblk2.b5_oRB_C[53]  (.D(mdiclink_reg[323]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[53]));
    SLE \genblk2.b5_oRB_C[64]  (.D(mdiclink_reg[312]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[64]));
    SLE \genblk2.b5_oRB_C[302]  (.D(mdiclink_reg[74]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[302]));
    SLE \genblk2.b5_oRB_C[293]  (.D(mdiclink_reg[83]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[293]));
    SLE \genblk2.b5_oRB_C[228]  (.D(mdiclink_reg[148]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[228]));
    SLE \genblk2.b5_oRB_C[116]  (.D(mdiclink_reg[260]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[116]));
    SLE \genblk2.b5_oRB_C[49]  (.D(mdiclink_reg[327]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[49]));
    SLE \genblk2.b5_oRB_C[99]  (.D(mdiclink_reg[277]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[99]));
    SLE \genblk2.b5_oRB_C[202]  (.D(mdiclink_reg[174]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[202]));
    VCC VCC (.Y(VCC_net_1));
    SLE \genblk2.b5_oRB_C[100]  (.D(mdiclink_reg[276]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[100]));
    SLE \genblk2.b5_oRB_C[279]  (.D(mdiclink_reg[97]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[279]));
    SLE \genblk2.b5_oRB_C[103]  (.D(mdiclink_reg[273]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[103]));
    SLE \genblk2.b5_oRB_C[156]  (.D(mdiclink_reg[220]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[156]));
    SLE \genblk2.b5_oRB_C[145]  (.D(mdiclink_reg[231]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[145]));
    SLE \genblk2.b5_oRB_C[55]  (.D(mdiclink_reg[321]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[55]));
    SLE \genblk2.b5_oRB_C[239]  (.D(mdiclink_reg[137]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[239]));
    SLE \genblk2.b5_oRB_C[364]  (.D(mdiclink_reg[12]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[364]));
    SLE \genblk2.b5_oRB_C[346]  (.D(mdiclink_reg[30]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[346]));
    SLE \genblk2.b5_oRB_C[194]  (.D(mdiclink_reg[182]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[194]));
    SLE \genblk2.b5_oRB_C[162]  (.D(mdiclink_reg[214]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[162]));
    SLE \genblk2.b5_oRB_C[309]  (.D(mdiclink_reg[67]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[309]));
    SLE \genblk2.b5_oRB_C[245]  (.D(mdiclink_reg[131]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[245]));
    SLE \genblk2.b5_oRB_C[27]  (.D(mdiclink_reg[349]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[27]));
    SLE \genblk2.b5_oRB_C[367]  (.D(mdiclink_reg[9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[367]));
    SLE \genblk2.b5_oRB_C[28]  (.D(mdiclink_reg[348]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[28]));
    SLE \genblk2.b5_oRB_C[14]  (.D(mdiclink_reg[362]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[14]));
    SLE \genblk2.b5_oRB_C[373]  (.D(mdiclink_reg[3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[373]));
    SLE \genblk2.b5_oRB_C[280]  (.D(mdiclink_reg[96]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[280]));
    SLE \genblk2.b5_oRB_C[333]  (.D(mdiclink_reg[43]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[333]));
    SLE \genblk2.b5_oRB_C[229]  (.D(mdiclink_reg[147]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[229]));
    SLE \genblk2.b5_oRB_C[368]  (.D(mdiclink_reg[8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[368]));
    SLE \genblk2.b5_oRB_C[266]  (.D(mdiclink_reg[110]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[266]));
    SLE \genblk2.b5_oRB_C[243]  (.D(mdiclink_reg[133]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[243]));
    SLE \genblk2.b5_oRB_C[37]  (.D(mdiclink_reg[339]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[37]));
    SLE \genblk2.b5_oRB_C[284]  (.D(mdiclink_reg[92]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[284]));
    SLE \genblk2.b5_oRB_C[196]  (.D(mdiclink_reg[180]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[196]));
    SLE \genblk2.b5_oRB_C[161]  (.D(mdiclink_reg[215]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[161]));
    SLE \genblk2.b5_oRB_C[188]  (.D(mdiclink_reg[188]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[188]));
    SLE \genblk2.b5_oRB_C[38]  (.D(mdiclink_reg[338]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[38]));
    SLE \genblk2.b5_oRB_C[69]  (.D(mdiclink_reg[307]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[69]));
    SLE \genblk2.b5_oRB_C[109]  (.D(mdiclink_reg[267]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[109]));
    SLE \genblk2.b5_oRB_C[1]  (.D(mdiclink_reg[375]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[1]));
    SLE \genblk2.b5_oRB_C[323]  (.D(mdiclink_reg[53]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[323]));
    SLE \genblk2.b5_oRB_C[210]  (.D(mdiclink_reg[166]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[210]));
    SLE \genblk2.b5_oRB_C[21]  (.D(mdiclink_reg[355]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[21]));
    SLE \genblk2.b5_oRB_C[167]  (.D(mdiclink_reg[209]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[167]));
    SLE \genblk2.b5_oRB_C[77]  (.D(mdiclink_reg[299]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[77]));
    SLE \genblk2.b5_oRB_C[144]  (.D(mdiclink_reg[232]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[144]));
    SLE \genblk2.b5_oRB_C[78]  (.D(mdiclink_reg[298]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[78]));
    SLE \genblk2.b5_oRB_C[87]  (.D(mdiclink_reg[289]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[87]));
    SLE \genblk2.b5_oRB_C[88]  (.D(mdiclink_reg[288]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[88]));
    SLE \genblk2.b5_oRB_C[42]  (.D(mdiclink_reg[334]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[42]));
    SLE \genblk2.b5_oRB_C[214]  (.D(mdiclink_reg[162]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[214]));
    SLE \genblk2.b5_oRB_C[92]  (.D(mdiclink_reg[284]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[92]));
    SLE \genblk2.b5_oRB_C[250]  (.D(mdiclink_reg[126]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[250]));
    SLE \genblk2.b5_oRB_C[118]  (.D(mdiclink_reg[258]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[118]));
    SLE \genblk2.b5_oRB_C[282]  (.D(mdiclink_reg[94]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[282]));
    SLE \genblk2.b5_oRB_C[26]  (.D(mdiclink_reg[350]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[26]));
    SLE \genblk2.b5_oRB_C[180]  (.D(mdiclink_reg[196]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[180]));
    SLE \genblk2.b5_oRB_C[31]  (.D(mdiclink_reg[345]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[31]));
    SLE \genblk2.b5_oRB_C[183]  (.D(mdiclink_reg[193]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[183]));
    SLE \genblk2.b5_oRB_C[315]  (.D(mdiclink_reg[61]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[315]));
    SLE \genblk2.b5_oRB_C[277]  (.D(mdiclink_reg[99]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[277]));
    SLE \genblk2.b5_oRB_C[254]  (.D(mdiclink_reg[122]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[254]));
    SLE \genblk2.b5_oRB_C[158]  (.D(mdiclink_reg[218]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[158]));
    SLE \genblk2.b5_oRB_C[237]  (.D(mdiclink_reg[139]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[237]));
    SLE \genblk2.b5_oRB_C[312]  (.D(mdiclink_reg[64]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[312]));
    SLE \genblk2.b5_oRB_C[36]  (.D(mdiclink_reg[340]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[36]));
    SLE \genblk2.b5_oRB_C[304]  (.D(mdiclink_reg[72]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[304]));
    SLE \genblk2.b5_oRB_C[146]  (.D(mdiclink_reg[230]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[146]));
    SLE \genblk2.b5_oRB_C[19]  (.D(mdiclink_reg[357]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[19]));
    SLE \genblk2.b5_oRB_C[9]  (.D(mdiclink_reg[367]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[9]));
    SLE \genblk2.b5_oRB_C[360]  (.D(mdiclink_reg[16]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[360]));
    SLE \genblk2.b5_oRB_C[71]  (.D(mdiclink_reg[305]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[71]));
    SLE \genblk2.b5_oRB_C[355]  (.D(mdiclink_reg[21]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[355]));
    SLE \genblk2.b5_oRB_C[102]  (.D(mdiclink_reg[274]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[102]));
    SLE \genblk2.b5_oRB_C[54]  (.D(mdiclink_reg[322]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[54]));
    SLE \genblk2.b5_oRB_C[81]  (.D(mdiclink_reg[295]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[81]));
    SLE \genblk2.b5_oRB_C[352]  (.D(mdiclink_reg[24]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[352]));
    SLE \genblk2.b5_oRB_C[212]  (.D(mdiclink_reg[164]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[212]));
    SLE \genblk2.b5_oRB_C[110]  (.D(mdiclink_reg[266]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[110]));
    SLE \genblk2.b5_oRB_C[307]  (.D(mdiclink_reg[69]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[307]));
    SLE \genblk2.b5_oRB_C[290]  (.D(mdiclink_reg[86]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[290]));
    SLE \genblk2.b5_oRB_C[113]  (.D(mdiclink_reg[263]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[113]));
    SLE \genblk2.b5_oRB_C[76]  (.D(mdiclink_reg[300]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[76]));
    SLE \genblk2.b5_oRB_C[227]  (.D(mdiclink_reg[149]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[227]));
    SLE \genblk2.b5_oRB_C[308]  (.D(mdiclink_reg[68]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[308]));
    SLE \genblk2.b5_oRB_C[86]  (.D(mdiclink_reg[290]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[86]));
    SLE \genblk2.b5_oRB_C[252]  (.D(mdiclink_reg[124]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[252]));
    SLE \genblk2.b5_oRB_C[206]  (.D(mdiclink_reg[170]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[206]));
    SLE \genblk2.b5_oRB_C[150]  (.D(mdiclink_reg[226]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[150]));
    SLE \genblk2.b5_oRB_C[294]  (.D(mdiclink_reg[82]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[294]));
    SLE \genblk2.b5_oRB_C[198]  (.D(mdiclink_reg[178]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[198]));
    SLE \genblk2.b5_oRB_C[175]  (.D(mdiclink_reg[201]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[175]));
    SLE \genblk2.b5_oRB_C[153]  (.D(mdiclink_reg[223]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[153]));
    SLE \genblk2.b5_oRB_C[101]  (.D(mdiclink_reg[275]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[101]));
    SLE \genblk2.b5_oRB_C[62]  (.D(mdiclink_reg[314]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[62]));
    SLE \genblk2.b5_oRB_C[319]  (.D(mdiclink_reg[57]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[319]));
    SLE \genblk2.b5_oRB_C[189]  (.D(mdiclink_reg[187]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[189]));
    SLE \genblk2.b5_oRB_C[135]  (.D(mdiclink_reg[241]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[135]));
    SLE \genblk2.b13_oRB_MqCD2_EdR  (.D(b13_oRB_MqCD2_EdR), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_2o_z));
    SLE \genblk2.b5_oRB_C[376]  (.D(mdiclink_reg[0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[376]));
    SLE \genblk2.b5_oRB_C[336]  (.D(mdiclink_reg[40]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[336]));
    SLE \genblk2.b5_oRB_C[275]  (.D(mdiclink_reg[101]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[275]));
    SLE \genblk2.b5_oRB_C[359]  (.D(mdiclink_reg[17]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[359]));
    SLE \genblk2.b5_oRB_C[235]  (.D(mdiclink_reg[141]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[235]));
    SLE \genblk2.b5_oRB_C[40]  (.D(mdiclink_reg[336]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[40]));
    SLE \genblk2.b5_oRB_C[107]  (.D(mdiclink_reg[269]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[107]));
    SLE \genblk2.b5_oRB_C[90]  (.D(mdiclink_reg[286]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[90]));
    SLE \genblk2.b5_oRB_C[23]  (.D(mdiclink_reg[353]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[23]));
    SLE \genblk2.b5_oRB_C[125]  (.D(mdiclink_reg[251]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[125]));
    SLE \genblk2.b5_oRB_C[292]  (.D(mdiclink_reg[84]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[292]));
    SLE \genblk2.b5_oRB_C[273]  (.D(mdiclink_reg[103]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[273]));
    SLE \genblk2.b5_oRB_C[190]  (.D(mdiclink_reg[186]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[190]));
    SLE \genblk2.b5_oRB_C[119]  (.D(mdiclink_reg[257]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[119]));
    SLE \genblk2.b5_oRB_C[326]  (.D(mdiclink_reg[50]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[326]));
    SLE \genblk2.b5_oRB_C[233]  (.D(mdiclink_reg[143]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[233]));
    SLE \genblk2.b5_oRB_C[240]  (.D(mdiclink_reg[136]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[240]));
    SLE \genblk2.b5_oRB_C[193]  (.D(mdiclink_reg[183]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[193]));
    SLE \genblk2.b5_oRB_C[33]  (.D(mdiclink_reg[343]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[33]));
    SLE \genblk2.b5_oRB_C[225]  (.D(mdiclink_reg[151]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[225]));
    SLE \genblk2.b5_oRB_C[59]  (.D(mdiclink_reg[317]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[59]));
    SLE \genblk2.b5_oRB_C[12]  (.D(mdiclink_reg[364]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[12]));
    SLE \genblk2.b5_oRB_C[361]  (.D(mdiclink_reg[15]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[361]));
    SLE \genblk2.b5_oRB_C[159]  (.D(mdiclink_reg[217]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[159]));
    SLE \genblk2.b5_oRB_C[244]  (.D(mdiclink_reg[132]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[244]));
    SLE \genblk2.b5_oRB_C[7]  (.D(mdiclink_reg[369]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[7]));
    SLE \genblk2.b5_oRB_C[25]  (.D(mdiclink_reg[351]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[25]));
    SLE \genblk2.b5_oRB_C[148]  (.D(mdiclink_reg[228]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[148]));
    SLE \genblk2.b5_oRB_C[261]  (.D(mdiclink_reg[115]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[261]));
    SLE \genblk2.b5_oRB_C[182]  (.D(mdiclink_reg[194]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[182]));
    SLE \genblk2.b5_oRB_C[300]  (.D(mdiclink_reg[76]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[300]));
    SLE \genblk2.b5_oRB_C[174]  (.D(mdiclink_reg[202]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[174]));
    SLE \genblk2.b5_oRB_C[223]  (.D(mdiclink_reg[153]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[223]));
    SLE \genblk2.b5_oRB_C[134]  (.D(mdiclink_reg[242]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[134]));
    SLE \genblk2.b5_oRB_C[73]  (.D(mdiclink_reg[303]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[73]));
    SLE \genblk2.b5_oRB_C[345]  (.D(mdiclink_reg[31]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[345]));
    SLE \genblk2.b5_oRB_C[83]  (.D(mdiclink_reg[293]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[83]));
    SLE \genblk2.b5_oRB_C[35]  (.D(mdiclink_reg[341]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[35]));
    SLE \genblk2.b5_oRB_C[342]  (.D(mdiclink_reg[34]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[342]));
    SLE \genblk2.b5_oRB_C[286]  (.D(mdiclink_reg[90]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[286]));
    SLE \genblk2.b5_oRB_C[60]  (.D(mdiclink_reg[316]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[60]));
    SLE \genblk2.b5_oRB_C[314]  (.D(mdiclink_reg[62]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[314]));
    SLE \genblk2.b5_oRB_C[181]  (.D(mdiclink_reg[195]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[181]));
    SLE \genblk2.b5_oRB_C[242]  (.D(mdiclink_reg[134]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[242]));
    SLE \genblk2.b5_oRB_C[112]  (.D(mdiclink_reg[264]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[112]));
    SLE \genblk2.b5_oRB_C[199]  (.D(mdiclink_reg[177]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[199]));
    SLE \genblk2.b5_oRB_C[140]  (.D(mdiclink_reg[236]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[140]));
    SLE \genblk2.b5_oRB_C[176]  (.D(mdiclink_reg[200]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[176]));
    SLE \genblk2.b5_oRB_C[143]  (.D(mdiclink_reg[233]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[143]));
    SLE \genblk2.b5_oRB_C[124]  (.D(mdiclink_reg[252]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[124]));
    SLE \genblk2.b5_oRB_C[75]  (.D(mdiclink_reg[301]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[75]));
    SLE \genblk2.b5_oRB_C[354]  (.D(mdiclink_reg[22]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[354]));
    SLE \genblk2.b5_oRB_C[317]  (.D(mdiclink_reg[59]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[317]));
    SLE \genblk2.b5_oRB_C[136]  (.D(mdiclink_reg[240]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[136]));
    SLE \genblk2.b5_oRB_C[85]  (.D(mdiclink_reg[291]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[85]));
    SLE \genblk2.b5_oRB_C[187]  (.D(mdiclink_reg[189]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[187]));
    SLE \genblk2.b5_oRB_C[152]  (.D(mdiclink_reg[224]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[152]));
    SLE \genblk2.b5_oRB_C[318]  (.D(mdiclink_reg[58]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[318]));
    SLE \genblk2.b5_oRB_C[216]  (.D(mdiclink_reg[160]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[216]));
    SLE \genblk2.b5_oRB_C[349]  (.D(mdiclink_reg[27]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[349]));
    SLE \genblk2.b5_oRB_C[357]  (.D(mdiclink_reg[19]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[357]));
    SLE \genblk2.b5_oRB_C[268]  (.D(mdiclink_reg[108]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[268]));
    SLE \genblk2.b5_oRB_C[111]  (.D(mdiclink_reg[265]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[111]));
    SLE \genblk2.b5_oRB_C[8]  (.D(mdiclink_reg[368]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[8]));
    SLE \genblk2.b5_oRB_C[358]  (.D(mdiclink_reg[18]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[358]));
    SLE \genblk2.b5_oRB_C[256]  (.D(mdiclink_reg[120]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[256]));
    SLE \genblk2.b5_oRB_C[2]  (.D(mdiclink_reg[374]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[2]));
    SLE \genblk2.b5_oRB_C[126]  (.D(mdiclink_reg[250]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[126]));
    SLE \genblk2.b5_oRB_C[10]  (.D(mdiclink_reg[366]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[10]));
    SLE \genblk2.b5_oRB_C[52]  (.D(mdiclink_reg[324]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[52]));
    SLE \genblk2.b5_oRB_C[151]  (.D(mdiclink_reg[225]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[151]));
    SLE \genblk2.b5_oRB_C[117]  (.D(mdiclink_reg[259]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[117]));
    SLE \genblk2.b5_oRB_C[301]  (.D(mdiclink_reg[75]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[301]));
    SLE \genblk2.b5_oRB_C[192]  (.D(mdiclink_reg[184]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[192]));
    SLE \genblk2.b5_oRB_C[201]  (.D(mdiclink_reg[175]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[201]));
    SLE \genblk2.b5_oRB_C[149]  (.D(mdiclink_reg[227]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[149]));
    SLE \genblk2.b5_oRB_C[157]  (.D(mdiclink_reg[219]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[157]));
    SLE \genblk2.b5_oRB_C[24]  (.D(mdiclink_reg[352]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[24]));
    CFG2 #( .INIT(4'hE) )  \genblk2.b13_oRB_MqCD2_EdR_s  (.A(
        b6_Ocm0rW_0_0_o2[2]), .B(b13_nAzGfFM_sLsv3[1]), .Y(
        b13_oRB_MqCD2_EdR));
    SLE \genblk2.b5_oRB_C[269]  (.D(mdiclink_reg[107]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[269]));
    SLE \genblk2.b5_oRB_C[296]  (.D(mdiclink_reg[80]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[296]));
    SLE \genblk2.b5_oRB_C[270]  (.D(mdiclink_reg[106]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[270]));
    SLE \genblk2.b5_oRB_C[191]  (.D(mdiclink_reg[185]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[191]));
    SLE \genblk2.b5_oRB_C[230]  (.D(mdiclink_reg[146]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[230]));
    SLE \genblk2.b5_oRB_C[310]  (.D(mdiclink_reg[66]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[310]));
    SLE \genblk2.b5_oRB_C[34]  (.D(mdiclink_reg[342]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[34]));
    SLE \genblk2.b5_oRB_C[274]  (.D(mdiclink_reg[102]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[274]));
    SLE \genblk2.b5_oRB_C[178]  (.D(mdiclink_reg[198]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[178]));
    SLE \genblk2.b5_oRB_C[234]  (.D(mdiclink_reg[142]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[234]));
    SLE \genblk2.b5_oRB_C[4]  (.D(mdiclink_reg[372]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[4]));
    SLE \genblk2.b5_oRB_C[138]  (.D(mdiclink_reg[238]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[138]));
    SLE \genblk2.b5_oRB_C[363]  (.D(mdiclink_reg[13]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[363]));
    SLE \genblk2.b5_oRB_C[350]  (.D(mdiclink_reg[26]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[350]));
    SLE \genblk2.b5_oRB_C[344]  (.D(mdiclink_reg[32]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[344]));
    SLE \genblk2.b5_oRB_C[197]  (.D(mdiclink_reg[179]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[197]));
    SLE \genblk2.b5_oRB_C[375]  (.D(mdiclink_reg[1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[375]));
    SLE \genblk2.b5_oRB_C[142]  (.D(mdiclink_reg[234]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[142]));
    SLE \genblk2.b5_oRB_C[74]  (.D(mdiclink_reg[302]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[74]));
    SLE \genblk2.b5_oRB_C[335]  (.D(mdiclink_reg[41]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[335]));
    SLE \genblk2.b5_oRB_C[220]  (.D(mdiclink_reg[156]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[220]));
    SLE \genblk2.b5_oRB_C[372]  (.D(mdiclink_reg[4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[372]));
    SLE \genblk2.b5_oRB_C[208]  (.D(mdiclink_reg[168]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[208]));
    SLE \genblk2.b5_oRB_C[84]  (.D(mdiclink_reg[292]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[84]));
    SLE \genblk2.b5_oRB_C[332]  (.D(mdiclink_reg[44]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[332]));
    SLE \genblk2.b5_oRB_C[50]  (.D(mdiclink_reg[326]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[50]));
    SLE \genblk2.b5_oRB_C[347]  (.D(mdiclink_reg[29]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[347]));
    SLE \genblk2.b5_oRB_C[224]  (.D(mdiclink_reg[152]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[224]));
    SLE \genblk2.b5_oRB_C[128]  (.D(mdiclink_reg[248]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[128]));
    SLE \genblk2.b5_oRB_C[348]  (.D(mdiclink_reg[28]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[348]));
    SLE \genblk2.b5_oRB_C[272]  (.D(mdiclink_reg[104]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[272]));
    SLE \genblk2.b5_oRB_C[246]  (.D(mdiclink_reg[130]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[246]));
    SLE \genblk2.b5_oRB_C[170]  (.D(mdiclink_reg[206]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[170]));
    SLE \genblk2.b5_oRB_C[232]  (.D(mdiclink_reg[144]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[232]));
    SLE \genblk2.b5_oRB_C[173]  (.D(mdiclink_reg[203]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[173]));
    SLE \genblk2.b5_oRB_C[130]  (.D(mdiclink_reg[246]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[130]));
    SLE \genblk2.b5_oRB_C[141]  (.D(mdiclink_reg[235]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[141]));
    SLE \genblk2.b5_oRB_C[133]  (.D(mdiclink_reg[243]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[133]));
    SLE \genblk2.b5_oRB_C[325]  (.D(mdiclink_reg[51]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[325]));
    SLE \genblk2.b5_oRB_C[281]  (.D(mdiclink_reg[95]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[281]));
    SLE \genblk2.b5_oRB_C[29]  (.D(mdiclink_reg[347]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[29]));
    SLE \genblk2.b5_oRB_C[322]  (.D(mdiclink_reg[54]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[322]));
    SLE \genblk2.b5_oRB_C[339]  (.D(mdiclink_reg[37]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[339]));
    SLE \genblk2.b5_oRB_C[147]  (.D(mdiclink_reg[229]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[147]));
    SLE \genblk2.b5_oRB_C[39]  (.D(mdiclink_reg[337]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[39]));
    SLE \genblk2.b5_oRB_C[222]  (.D(mdiclink_reg[154]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[222]));
    SLE \genblk2.b5_oRB_C[267]  (.D(mdiclink_reg[109]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[267]));
    SLE \genblk2.b5_oRB_C[209]  (.D(mdiclink_reg[167]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[209]));
    SLE \genblk2.b5_oRB_C[120]  (.D(mdiclink_reg[256]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[120]));
    SLE \genblk2.b5_oRB_C[311]  (.D(mdiclink_reg[65]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[311]));
    SLE \genblk2.b5_oRB_C[123]  (.D(mdiclink_reg[253]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[123]));
    SLE \genblk2.b5_oRB_C[47]  (.D(mdiclink_reg[329]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[47]));
    SLE \genblk2.b5_oRB_C[97]  (.D(mdiclink_reg[279]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[97]));
    SLE \genblk2.b5_oRB_C[211]  (.D(mdiclink_reg[165]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[211]));
    SLE \genblk2.b5_oRB_C[48]  (.D(mdiclink_reg[328]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[48]));
    SLE \genblk2.b5_oRB_C[98]  (.D(mdiclink_reg[278]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[98]));
    SLE \genblk2.b5_oRB_C[351]  (.D(mdiclink_reg[25]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[351]));
    SLE \genblk2.b5_oRB_C[79]  (.D(mdiclink_reg[297]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[79]));
    SLE \genblk2.b5_oRB_C[329]  (.D(mdiclink_reg[47]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[329]));
    SLE \genblk2.b5_oRB_C[179]  (.D(mdiclink_reg[197]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[179]));
    SLE \genblk2.b5_oRB_C[251]  (.D(mdiclink_reg[125]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[251]));
    SLE \genblk2.b5_oRB_C[89]  (.D(mdiclink_reg[287]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[89]));
    SLE \genblk2.b5_oRB_C[139]  (.D(mdiclink_reg[237]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[139]));
    SLE \genblk2.b5_oRB_C[303]  (.D(mdiclink_reg[73]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[303]));
    SLE \genblk2.b5_oRB_C[340]  (.D(mdiclink_reg[36]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[340]));
    SLE \genblk2.b5_oRB_C[288]  (.D(mdiclink_reg[88]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[288]));
    SLE \genblk2.b5_oRB_C[165]  (.D(mdiclink_reg[211]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[165]));
    SLE \genblk2.b5_oRB_C[6]  (.D(mdiclink_reg[370]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[6]));
    SLE \genblk2.b5_oRB_C[41]  (.D(mdiclink_reg[335]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[41]));
    SLE \genblk2.b5_oRB_C[366]  (.D(mdiclink_reg[10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[366]));
    SLE \genblk2.b5_oRB_C[91]  (.D(mdiclink_reg[285]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[91]));
    SLE \genblk2.b5_oRB_C[129]  (.D(mdiclink_reg[247]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[129]));
    SLE \genblk2.b5_oRB_C[265]  (.D(mdiclink_reg[111]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[265]));
    SLE \genblk2.b5_oRB_C[22]  (.D(mdiclink_reg[354]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[22]));
    SLE \genblk2.b5_oRB_C[46]  (.D(mdiclink_reg[330]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[46]));
    SLE \genblk2.b5_oRB_C[96]  (.D(mdiclink_reg[280]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[96]));
    SLE \genblk2.b5_oRB_C[291]  (.D(mdiclink_reg[85]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[291]));
    SLE \genblk2.b5_oRB_C[67]  (.D(mdiclink_reg[309]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[67]));
    SLE \genblk2.b5_oRB_C[374]  (.D(mdiclink_reg[2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[374]));
    SLE \genblk2.b5_oRB_C[218]  (.D(mdiclink_reg[158]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[218]));
    SLE \genblk2.b5_oRB_C[68]  (.D(mdiclink_reg[308]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[68]));
    SLE \genblk2.b5_oRB_C[334]  (.D(mdiclink_reg[42]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[334]));
    SLE \genblk2.b5_oRB_C[263]  (.D(mdiclink_reg[113]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[263]));
    SLE \genblk2.b5_oRB_C[172]  (.D(mdiclink_reg[204]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[172]));
    SLE \genblk2.b5_oRB_C[32]  (.D(mdiclink_reg[344]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[32]));
    SLE \genblk2.b5_oRB_C[132]  (.D(mdiclink_reg[244]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[132]));
    SLE \genblk2.b5_oRB_C[289]  (.D(mdiclink_reg[87]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[289]));
    SLE \genblk2.b5_oRB_C[258]  (.D(mdiclink_reg[118]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[258]));
    
endmodule


module b11_OFWNT9s_8tZ_Z2_x(
       b11_OFWNT9L_8tZ,
       mdiclink_reg,
       b6_Ocm0rW_0_0_o2,
       b13_nAzGfFM_sLsv3,
       IICE_comm2iice_11,
       IICE_comm2iice_10,
       IICE_comm2iice_5,
       IICE_comm2iice_0,
       IICE_comm2iice_4,
       IICE_comm2iice_9,
       IICE_comm2iice_1,
       IICE_comm2iice_3,
       IICE_comm2iice_2,
       IICE_comm2iice_6,
       BW_clk_c,
       b11_PSyil9s_FMZ,
       b8_SoWGfWYY_i,
       b8_SoWGfWYY,
       b10_OFWNT9khFt,
       b7_yYh03wy,
       b9_OFWNT9Mxf
    );
output [376:0] b11_OFWNT9L_8tZ;
input  [376:0] mdiclink_reg;
input  [2:2] b6_Ocm0rW_0_0_o2;
input  [1:1] b13_nAzGfFM_sLsv3;
input  IICE_comm2iice_11;
input  IICE_comm2iice_10;
input  IICE_comm2iice_5;
input  IICE_comm2iice_0;
input  IICE_comm2iice_4;
input  IICE_comm2iice_9;
input  IICE_comm2iice_1;
input  IICE_comm2iice_3;
input  IICE_comm2iice_2;
input  IICE_comm2iice_6;
input  BW_clk_c;
input  b11_PSyil9s_FMZ;
input  b8_SoWGfWYY_i;
input  b8_SoWGfWYY;
input  b10_OFWNT9khFt;
output b7_yYh03wy;
output b9_OFWNT9Mxf;

    wire \b12_PSyi_KyDbLbb[0]_net_1 , VCC_net_1, 
        \b12_2_St6KCa_jHv[0]_net_1 , b12_PSyi_KyDbLbb_0_sqmuxa_net_1, 
        GND_net_1, \b12_PSyi_KyDbLbb[1]_net_1 , 
        \b12_2_St6KCa_jHv[1]_net_1 , \b12_PSyi_KyDbLbb[2]_net_1 , 
        \b12_2_St6KCa_jHv[2]_net_1 , \b12_PSyi_KyDbLbb[3]_net_1 , 
        \b12_2_St6KCa_jHv[3]_net_1 , \b12_PSyi_KyDbLbb[4]_net_1 , 
        \b12_2_St6KCa_jHv[4]_net_1 , \b12_PSyi_KyDbLbb[5]_net_1 , 
        \b12_2_St6KCa_jHv[5]_net_1 , \b12_PSyi_KyDbLbb[6]_net_1 , 
        \b12_2_St6KCa_jHv[6]_net_1 , \b12_PSyi_KyDbLbb[7]_net_1 , 
        \b12_2_St6KCa_jHv[7]_net_1 , \b12_PSyi_KyDbLbb[8]_net_1 , 
        \b12_2_St6KCa_jHv[8]_net_1 , \b12_PSyi_KyDbLbb[9]_net_1 , 
        \b12_2_St6KCa_jHv[9]_net_1 , b9_PSyil9s_2_net_1, b8_nYJ_TqLY, 
        \b7_nYJ_BFM[382] , \b7_nYJ_BFM_or[7] , \b7_nYJ_BFM[368] , 
        \b7_nYJ_BFM[367] , \b7_nYJ_BFM[369] , \b7_nYJ_BFM[370] , 
        \b7_nYJ_BFM[371] , \b7_nYJ_BFM[372] , \b7_nYJ_BFM[373] , 
        \b7_nYJ_BFM[374] , \b7_nYJ_BFM[375] , \b7_nYJ_BFM[376] , 
        \b7_nYJ_BFM[377] , \b7_nYJ_BFM[378] , \b7_nYJ_BFM[379] , 
        \b7_nYJ_BFM[380] , \b7_nYJ_BFM[381] , \b7_nYJ_BFM[353] , 
        \b7_nYJ_BFM[352] , \b7_nYJ_BFM[354] , \b7_nYJ_BFM[355] , 
        \b7_nYJ_BFM[356] , \b7_nYJ_BFM[357] , \b7_nYJ_BFM[358] , 
        \b7_nYJ_BFM[359] , \b7_nYJ_BFM[360] , \b7_nYJ_BFM[361] , 
        \b7_nYJ_BFM[362] , \b7_nYJ_BFM[363] , \b7_nYJ_BFM[364] , 
        \b7_nYJ_BFM[365] , \b7_nYJ_BFM[366] , \b7_nYJ_BFM[338] , 
        \b7_nYJ_BFM[337] , \b7_nYJ_BFM[339] , \b7_nYJ_BFM[340] , 
        \b7_nYJ_BFM[341] , \b7_nYJ_BFM[342] , \b7_nYJ_BFM[343] , 
        \b7_nYJ_BFM[344] , \b7_nYJ_BFM[345] , \b7_nYJ_BFM[346] , 
        \b7_nYJ_BFM[347] , \b7_nYJ_BFM[348] , \b7_nYJ_BFM[349] , 
        \b7_nYJ_BFM[350] , \b7_nYJ_BFM[351] , \b7_nYJ_BFM[323] , 
        \b7_nYJ_BFM[322] , \b7_nYJ_BFM[324] , \b7_nYJ_BFM[325] , 
        \b7_nYJ_BFM[326] , \b7_nYJ_BFM[327] , \b7_nYJ_BFM[328] , 
        \b7_nYJ_BFM[329] , \b7_nYJ_BFM[330] , \b7_nYJ_BFM[331] , 
        \b7_nYJ_BFM[332] , \b7_nYJ_BFM[333] , \b7_nYJ_BFM[334] , 
        \b7_nYJ_BFM[335] , \b7_nYJ_BFM[336] , \b7_nYJ_BFM[308] , 
        \b7_nYJ_BFM[307] , \b7_nYJ_BFM[309] , \b7_nYJ_BFM[310] , 
        \b7_nYJ_BFM[311] , \b7_nYJ_BFM[312] , \b7_nYJ_BFM[313] , 
        \b7_nYJ_BFM[314] , \b7_nYJ_BFM[315] , \b7_nYJ_BFM[316] , 
        \b7_nYJ_BFM[317] , \b7_nYJ_BFM[318] , \b7_nYJ_BFM[319] , 
        \b7_nYJ_BFM[320] , \b7_nYJ_BFM[321] , \b7_nYJ_BFM[293] , 
        \b7_nYJ_BFM[292] , \b7_nYJ_BFM[294] , \b7_nYJ_BFM[295] , 
        \b7_nYJ_BFM[296] , \b7_nYJ_BFM[297] , \b7_nYJ_BFM[298] , 
        \b7_nYJ_BFM[299] , \b7_nYJ_BFM[300] , \b7_nYJ_BFM[301] , 
        \b7_nYJ_BFM[302] , \b7_nYJ_BFM[303] , \b7_nYJ_BFM[304] , 
        \b7_nYJ_BFM[305] , \b7_nYJ_BFM[306] , \b7_nYJ_BFM[278] , 
        \b7_nYJ_BFM[277] , \b7_nYJ_BFM[279] , \b7_nYJ_BFM[280] , 
        \b7_nYJ_BFM[281] , \b7_nYJ_BFM[282] , \b7_nYJ_BFM[283] , 
        \b7_nYJ_BFM[284] , \b7_nYJ_BFM[285] , \b7_nYJ_BFM[286] , 
        \b7_nYJ_BFM[287] , \b7_nYJ_BFM[288] , \b7_nYJ_BFM[289] , 
        \b7_nYJ_BFM[290] , \b7_nYJ_BFM[291] , \b7_nYJ_BFM[263] , 
        \b7_nYJ_BFM[262] , \b7_nYJ_BFM[264] , \b7_nYJ_BFM[265] , 
        \b7_nYJ_BFM[266] , \b7_nYJ_BFM[267] , \b7_nYJ_BFM[268] , 
        \b7_nYJ_BFM[269] , \b7_nYJ_BFM[270] , \b7_nYJ_BFM[271] , 
        \b7_nYJ_BFM[272] , \b7_nYJ_BFM[273] , \b7_nYJ_BFM[274] , 
        \b7_nYJ_BFM[275] , \b7_nYJ_BFM[276] , \b7_nYJ_BFM[248] , 
        \b7_nYJ_BFM[247] , \b7_nYJ_BFM[249] , \b7_nYJ_BFM[250] , 
        \b7_nYJ_BFM[251] , \b7_nYJ_BFM[252] , \b7_nYJ_BFM[253] , 
        \b7_nYJ_BFM[254] , \b7_nYJ_BFM[255] , \b7_nYJ_BFM[256] , 
        \b7_nYJ_BFM[257] , \b7_nYJ_BFM[258] , \b7_nYJ_BFM[259] , 
        \b7_nYJ_BFM[260] , \b7_nYJ_BFM[261] , \b7_nYJ_BFM[233] , 
        \b7_nYJ_BFM[232] , \b7_nYJ_BFM[234] , \b7_nYJ_BFM[235] , 
        \b7_nYJ_BFM[236] , \b7_nYJ_BFM[237] , \b7_nYJ_BFM[238] , 
        \b7_nYJ_BFM[239] , \b7_nYJ_BFM[240] , \b7_nYJ_BFM[241] , 
        \b7_nYJ_BFM[242] , \b7_nYJ_BFM[243] , \b7_nYJ_BFM[244] , 
        \b7_nYJ_BFM[245] , \b7_nYJ_BFM[246] , \b7_nYJ_BFM[218] , 
        \b7_nYJ_BFM[217] , \b7_nYJ_BFM[219] , \b7_nYJ_BFM[220] , 
        \b7_nYJ_BFM[221] , \b7_nYJ_BFM[222] , \b7_nYJ_BFM[223] , 
        \b7_nYJ_BFM[224] , \b7_nYJ_BFM[225] , \b7_nYJ_BFM[226] , 
        \b7_nYJ_BFM[227] , \b7_nYJ_BFM[228] , \b7_nYJ_BFM[229] , 
        \b7_nYJ_BFM[230] , \b7_nYJ_BFM[231] , \b7_nYJ_BFM[203] , 
        \b7_nYJ_BFM[202] , \b7_nYJ_BFM[204] , \b7_nYJ_BFM[205] , 
        \b7_nYJ_BFM[206] , \b7_nYJ_BFM[207] , \b7_nYJ_BFM[208] , 
        \b7_nYJ_BFM[209] , \b7_nYJ_BFM[210] , \b7_nYJ_BFM[211] , 
        \b7_nYJ_BFM[212] , \b7_nYJ_BFM[213] , \b7_nYJ_BFM[214] , 
        \b7_nYJ_BFM[215] , \b7_nYJ_BFM[216] , \b7_nYJ_BFM[188] , 
        \b7_nYJ_BFM[187] , \b7_nYJ_BFM[189] , \b7_nYJ_BFM[190] , 
        \b7_nYJ_BFM[191] , \b7_nYJ_BFM[192] , \b7_nYJ_BFM[193] , 
        \b7_nYJ_BFM[194] , \b7_nYJ_BFM[195] , \b7_nYJ_BFM[196] , 
        \b7_nYJ_BFM[197] , \b7_nYJ_BFM[198] , \b7_nYJ_BFM[199] , 
        \b7_nYJ_BFM[200] , \b7_nYJ_BFM[201] , \b7_nYJ_BFM[173] , 
        \b7_nYJ_BFM[172] , \b7_nYJ_BFM[174] , \b7_nYJ_BFM[175] , 
        \b7_nYJ_BFM[176] , \b7_nYJ_BFM[177] , \b7_nYJ_BFM[178] , 
        \b7_nYJ_BFM[179] , \b7_nYJ_BFM[180] , \b7_nYJ_BFM[181] , 
        \b7_nYJ_BFM[182] , \b7_nYJ_BFM[183] , \b7_nYJ_BFM[184] , 
        \b7_nYJ_BFM[185] , \b7_nYJ_BFM[186] , \b7_nYJ_BFM[158] , 
        \b7_nYJ_BFM[157] , \b7_nYJ_BFM[159] , \b7_nYJ_BFM[160] , 
        \b7_nYJ_BFM[161] , \b7_nYJ_BFM[162] , \b7_nYJ_BFM[163] , 
        \b7_nYJ_BFM[164] , \b7_nYJ_BFM[165] , \b7_nYJ_BFM[166] , 
        \b7_nYJ_BFM[167] , \b7_nYJ_BFM[168] , \b7_nYJ_BFM[169] , 
        \b7_nYJ_BFM[170] , \b7_nYJ_BFM[171] , \b7_nYJ_BFM[143] , 
        \b7_nYJ_BFM[142] , \b7_nYJ_BFM[144] , \b7_nYJ_BFM[145] , 
        \b7_nYJ_BFM[146] , \b7_nYJ_BFM[147] , \b7_nYJ_BFM[148] , 
        \b7_nYJ_BFM[149] , \b7_nYJ_BFM[150] , \b7_nYJ_BFM[151] , 
        \b7_nYJ_BFM[152] , \b7_nYJ_BFM[153] , \b7_nYJ_BFM[154] , 
        \b7_nYJ_BFM[155] , \b7_nYJ_BFM[156] , \b7_nYJ_BFM[128] , 
        \b7_nYJ_BFM[127] , \b7_nYJ_BFM[129] , \b7_nYJ_BFM[130] , 
        \b7_nYJ_BFM[131] , \b7_nYJ_BFM[132] , \b7_nYJ_BFM[133] , 
        \b7_nYJ_BFM[134] , \b7_nYJ_BFM[135] , \b7_nYJ_BFM[136] , 
        \b7_nYJ_BFM[137] , \b7_nYJ_BFM[138] , \b7_nYJ_BFM[139] , 
        \b7_nYJ_BFM[140] , \b7_nYJ_BFM[141] , \b7_nYJ_BFM[113] , 
        \b7_nYJ_BFM[112] , \b7_nYJ_BFM[114] , \b7_nYJ_BFM[115] , 
        \b7_nYJ_BFM[116] , \b7_nYJ_BFM[117] , \b7_nYJ_BFM[118] , 
        \b7_nYJ_BFM[119] , \b7_nYJ_BFM[120] , \b7_nYJ_BFM[121] , 
        \b7_nYJ_BFM[122] , \b7_nYJ_BFM[123] , \b7_nYJ_BFM[124] , 
        \b7_nYJ_BFM[125] , \b7_nYJ_BFM[126] , \b7_nYJ_BFM[98] , 
        \b7_nYJ_BFM[97] , \b7_nYJ_BFM[99] , \b7_nYJ_BFM[100] , 
        \b7_nYJ_BFM[101] , \b7_nYJ_BFM[102] , \b7_nYJ_BFM[103] , 
        \b7_nYJ_BFM[104] , \b7_nYJ_BFM[105] , \b7_nYJ_BFM[106] , 
        \b7_nYJ_BFM[107] , \b7_nYJ_BFM[108] , \b7_nYJ_BFM[109] , 
        \b7_nYJ_BFM[110] , \b7_nYJ_BFM[111] , \b7_nYJ_BFM[83] , 
        \b7_nYJ_BFM[82] , \b7_nYJ_BFM[84] , \b7_nYJ_BFM[85] , 
        \b7_nYJ_BFM[86] , \b7_nYJ_BFM[87] , \b7_nYJ_BFM[88] , 
        \b7_nYJ_BFM[89] , \b7_nYJ_BFM[90] , \b7_nYJ_BFM[91] , 
        \b7_nYJ_BFM[92] , \b7_nYJ_BFM[93] , \b7_nYJ_BFM[94] , 
        \b7_nYJ_BFM[95] , \b7_nYJ_BFM[96] , \b7_nYJ_BFM[68] , 
        \b7_nYJ_BFM[67] , \b7_nYJ_BFM[69] , \b7_nYJ_BFM[70] , 
        \b7_nYJ_BFM[71] , \b7_nYJ_BFM[72] , \b7_nYJ_BFM[73] , 
        \b7_nYJ_BFM[74] , \b7_nYJ_BFM[75] , \b7_nYJ_BFM[76] , 
        \b7_nYJ_BFM[77] , \b7_nYJ_BFM[78] , \b7_nYJ_BFM[79] , 
        \b7_nYJ_BFM[80] , \b7_nYJ_BFM[81] , \b7_nYJ_BFM[53] , 
        \b7_nYJ_BFM[52] , \b7_nYJ_BFM[54] , \b7_nYJ_BFM[55] , 
        \b7_nYJ_BFM[56] , \b7_nYJ_BFM[57] , \b7_nYJ_BFM[58] , 
        \b7_nYJ_BFM[59] , \b7_nYJ_BFM[60] , \b7_nYJ_BFM[61] , 
        \b7_nYJ_BFM[62] , \b7_nYJ_BFM[63] , \b7_nYJ_BFM[64] , 
        \b7_nYJ_BFM[65] , \b7_nYJ_BFM[66] , \b7_nYJ_BFM[38] , 
        \b7_nYJ_BFM[37] , \b7_nYJ_BFM[39] , \b7_nYJ_BFM[40] , 
        \b7_nYJ_BFM[41] , \b7_nYJ_BFM[42] , \b7_nYJ_BFM[43] , 
        \b7_nYJ_BFM[44] , \b7_nYJ_BFM[45] , \b7_nYJ_BFM[46] , 
        \b7_nYJ_BFM[47] , \b7_nYJ_BFM[48] , \b7_nYJ_BFM[49] , 
        \b7_nYJ_BFM[50] , \b7_nYJ_BFM[51] , \b7_nYJ_BFM[23] , 
        \b7_nYJ_BFM[22] , \b7_nYJ_BFM[24] , \b7_nYJ_BFM[25] , 
        \b7_nYJ_BFM[26] , \b7_nYJ_BFM[27] , \b7_nYJ_BFM[28] , 
        \b7_nYJ_BFM[29] , \b7_nYJ_BFM[30] , \b7_nYJ_BFM[31] , 
        \b7_nYJ_BFM[32] , \b7_nYJ_BFM[33] , \b7_nYJ_BFM[34] , 
        \b7_nYJ_BFM[35] , \b7_nYJ_BFM[36] , \b7_nYJ_BFM[8] , 
        \b7_nYJ_BFM[7] , \b7_nYJ_BFM[9] , \b7_nYJ_BFM[10] , 
        \b7_nYJ_BFM[11] , \b7_nYJ_BFM[12] , \b7_nYJ_BFM[13] , 
        \b7_nYJ_BFM[14] , \b7_nYJ_BFM[15] , \b7_nYJ_BFM[16] , 
        \b7_nYJ_BFM[17] , \b7_nYJ_BFM[18] , \b7_nYJ_BFM[19] , 
        \b7_nYJ_BFM[20] , \b7_nYJ_BFM[21] , \b8_FZFFLXYE[3]_net_1 , 
        b13_oRB_MqCD2_EdR_RNI9OIA, \b8_FZFFLXYE[4]_net_1 , 
        \b8_FZFFLXYE[5]_net_1 , \b8_FZFFLXYE[6]_net_1 , 
        \b8_FZFFLXYE[7]_net_1 , \b8_FZFFLXYE[8]_net_1 , 
        \b8_FZFFLXYE[9]_net_1 , \b7_nYJ_BFM[0] , \b7_nYJ_BFM[1] , 
        \b7_nYJ_BFM[2] , \b7_nYJ_BFM[3] , \b7_nYJ_BFM[4] , 
        \b7_nYJ_BFM[5] , \b7_nYJ_BFM[6] , N_850_a2_1_net_1, 
        \b8_FZFFLXYE[0]_net_1 , \b8_FZFFLXYE[1]_net_1 , 
        \b8_FZFFLXYE[2]_net_1 , b8_jAA_KlCO_net_1, 
        b8_jAA_KlCO_RNO_net_1, b8_jAA_KlCO_0_sqmuxa_net_1, 
        \b9_v_mzCDYXs[4] , b9_v_mzCDYXs_8, \b9_v_mzCDYXs[5] , 
        b9_v_mzCDYXs_7, \b9_v_mzCDYXs[6] , b9_v_mzCDYXs_6, 
        \b9_v_mzCDYXs[7] , b9_v_mzCDYXs_5, \b9_v_mzCDYXs[8] , 
        b9_v_mzCDYXs_4, \b9_v_mzCDYXs[9] , b9_v_mzCDYXs_3, 
        \b9_v_mzCDYXs[0] , b9_v_mzCDYXs_2, \b9_v_mzCDYXs[1] , 
        b9_v_mzCDYXs_1, \b9_v_mzCDYXs[2] , b9_v_mzCDYXs_0, 
        \b9_v_mzCDYXs[3] , b9_v_mzCDYXs, b12_2_St6KCa_jHv_8, 
        b12_2_St6KCa_jHv_7, b12_2_St6KCa_jHv_6, b12_2_St6KCa_jHv_5, 
        b12_2_St6KCa_jHv_4, b12_2_St6KCa_jHv_3, b12_2_St6KCa_jHv_2, 
        b12_2_St6KCa_jHv_1, b12_2_St6KCa_jHv_0, b12_2_St6KCa_jHv, 
        b9_v_mzCDYXs_cry_0_cy, N_24_mux, b9_v_mzCDYXs_cry_0, 
        \b9_v_mzCDYXs_RNIUDLP4_S[0] , b9_v_mzCDYXs_cry_1, 
        \b9_v_mzCDYXs_RNIA2R45_S[1] , b9_v_mzCDYXs_cry_2, 
        \b9_v_mzCDYXs_RNINN0G5_S[2] , b9_v_mzCDYXs_cry_3, 
        \b9_v_mzCDYXs_RNI5E6R5_S[3] , b9_v_mzCDYXs_cry_4, 
        \b9_v_mzCDYXs_RNIK5C66_S[4] , b9_v_mzCDYXs_cry_5, 
        \b9_v_mzCDYXs_RNI4UHH6_S[5] , b9_v_mzCDYXs_cry_6, 
        \b9_v_mzCDYXs_RNILNNS6_S[6] , b9_v_mzCDYXs_cry_7, 
        \b9_v_mzCDYXs_RNI7IT77_S[7] , \b9_v_mzCDYXs_r_RNO_S[9] , 
        b9_v_mzCDYXs_cry_8, \b9_v_mzCDYXs_RNIQD3J7_S[8] , 
        un1_b12_2_St6KCa_jHv_s_0_532_FCO, b4_2o_z, 
        un1_b12_2_St6KCa_jHv_cry_0_net_1, un1_b12_2_St6KCa_jHv_cry_0_S, 
        un1_b12_2_St6KCa_jHv_cry_1_net_1, un1_b12_2_St6KCa_jHv_cry_1_S, 
        un1_b12_2_St6KCa_jHv_cry_2_net_1, un1_b12_2_St6KCa_jHv_cry_2_S, 
        un1_b12_2_St6KCa_jHv_cry_3_net_1, un1_b12_2_St6KCa_jHv_cry_3_S, 
        un1_b12_2_St6KCa_jHv_cry_4_net_1, un1_b12_2_St6KCa_jHv_cry_4_S, 
        un1_b12_2_St6KCa_jHv_cry_5_net_1, un1_b12_2_St6KCa_jHv_cry_5_S, 
        un1_b12_2_St6KCa_jHv_cry_6_net_1, un1_b12_2_St6KCa_jHv_cry_6_S, 
        un1_b12_2_St6KCa_jHv_cry_7_net_1, un1_b12_2_St6KCa_jHv_cry_7_S, 
        un1_b12_2_St6KCa_jHv_s_9_S, un1_b12_2_St6KCa_jHv_cry_8_net_1, 
        un1_b12_2_St6KCa_jHv_cry_8_S, \b7_nYJ_BFM_RNI95U74[383] , 
        b8_jAA_KlCO_0_sqmuxa_4_net_1, \b7_vFW_PlM[265] , 
        \un1_b4_BVmQ[265] , \b7_vFW_PlM[1] , \un1_b4_BVmQ[1] , b4_ycsM, 
        ttdo, b7_yYh03wy_u_0_m2_net_1, \b7_vFW_PlM[263] , 
        \b7_vFW_PlM[7] , b3_PLF_187_net_1, \b7_vFW_PlM[136] , 
        \b7_vFW_PlM[9] , b3_PLF_186_net_1, \b7_vFW_PlM[282] , 
        \b7_vFW_PlM[171] , b3_PLF_184_net_1, \b7_vFW_PlM[316] , 
        \b7_vFW_PlM[60] , b3_PLF_183_net_1, \b7_vFW_PlM[205] , 
        \b7_vFW_PlM[94] , b3_PLF_182_net_1, \b7_vFW_PlM[350] , 
        \b7_vFW_PlM[239] , b3_PLF_181_net_1, \b7_vFW_PlM[368] , 
        \b7_vFW_PlM[112] , b3_PLF_180_net_1, \b7_vFW_PlM[241] , 
        \b7_vFW_PlM[114] , b3_PLF_179_net_1, \b7_vFW_PlM[370] , 
        \b7_vFW_PlM[243] , b3_PLF_178_net_1, \b7_vFW_PlM[372] , 
        \b7_vFW_PlM[116] , b3_PLF_177_net_1, \b7_vFW_PlM[245] , 
        \b7_vFW_PlM[118] , b3_PLF_176_net_1, \b7_vFW_PlM[374] , 
        \b7_vFW_PlM[247] , b3_PLF_175_net_1, \b7_vFW_PlM[376] , 
        \b7_vFW_PlM[120] , b3_PLF_174_net_1, \b7_vFW_PlM[249] , 
        \b7_vFW_PlM[138] , b3_PLF_173_net_1, \b7_vFW_PlM[155] , 
        \b7_vFW_PlM[44] , b3_PLF_172_net_1, \b7_vFW_PlM[300] , 
        \b7_vFW_PlM[189] , b3_PLF_171_net_1, \b7_vFW_PlM[334] , 
        \b7_vFW_PlM[78] , b3_PLF_170_net_1, \b7_vFW_PlM[223] , 
        \b7_vFW_PlM[96] , b3_PLF_169_net_1, \b7_vFW_PlM[352] , 
        \b7_vFW_PlM[225] , b3_PLF_168_net_1, \b7_vFW_PlM[354] , 
        \b7_vFW_PlM[98] , b3_PLF_167_net_1, \b7_vFW_PlM[227] , 
        \b7_vFW_PlM[100] , b3_PLF_166_net_1, \b7_vFW_PlM[356] , 
        \b7_vFW_PlM[229] , b3_PLF_165_net_1, \b7_vFW_PlM[358] , 
        \b7_vFW_PlM[102] , b3_PLF_164_net_1, \b7_vFW_PlM[231] , 
        \b7_vFW_PlM[104] , b3_PLF_163_net_1, \b7_vFW_PlM[360] , 
        \b7_vFW_PlM[233] , b3_PLF_162_net_1, \b7_vFW_PlM[139] , 
        \b7_vFW_PlM[122] , b3_PLF_161_net_1, \b7_vFW_PlM[284] , 
        \b7_vFW_PlM[28] , b3_PLF_160_net_1, \b7_vFW_PlM[173] , 
        \b7_vFW_PlM[62] , b3_PLF_159_net_1, \b7_vFW_PlM[318] , 
        \b7_vFW_PlM[207] , b3_PLF_158_net_1, \b7_vFW_PlM[336] , 
        \b7_vFW_PlM[80] , b3_PLF_157_net_1, \b7_vFW_PlM[209] , 
        \b7_vFW_PlM[82] , b3_PLF_156_net_1, \b7_vFW_PlM[338] , 
        \b7_vFW_PlM[211] , b3_PLF_155_net_1, \b7_vFW_PlM[340] , 
        \b7_vFW_PlM[84] , b3_PLF_154_net_1, \b7_vFW_PlM[213] , 
        \b7_vFW_PlM[86] , b3_PLF_153_net_1, \b7_vFW_PlM[342] , 
        \b7_vFW_PlM[215] , b3_PLF_152_net_1, \b7_vFW_PlM[344] , 
        \b7_vFW_PlM[88] , b3_PLF_151_net_1, \b7_vFW_PlM[217] , 
        \b7_vFW_PlM[106] , b3_PLF_150_net_1, \b7_vFW_PlM[363] , 
        \b7_vFW_PlM[123] , b3_PLF_149_net_1, \b7_vFW_PlM[268] , 
        \b7_vFW_PlM[157] , b3_PLF_148_net_1, \b7_vFW_PlM[302] , 
        \b7_vFW_PlM[46] , b3_PLF_147_net_1, \b7_vFW_PlM[191] , 
        \b7_vFW_PlM[64] , b3_PLF_146_net_1, \b7_vFW_PlM[320] , 
        \b7_vFW_PlM[193] , b3_PLF_145_net_1, \b7_vFW_PlM[322] , 
        \b7_vFW_PlM[66] , b3_PLF_144_net_1, \b7_vFW_PlM[195] , 
        \b7_vFW_PlM[68] , b3_PLF_143_net_1, \b7_vFW_PlM[324] , 
        \b7_vFW_PlM[197] , b3_PLF_142_net_1, \b7_vFW_PlM[326] , 
        \b7_vFW_PlM[70] , b3_PLF_141_net_1, \b7_vFW_PlM[199] , 
        \b7_vFW_PlM[72] , b3_PLF_140_net_1, \b7_vFW_PlM[328] , 
        \b7_vFW_PlM[201] , b3_PLF_139_net_1, \b7_vFW_PlM[107] , 
        \b7_vFW_PlM[90] , b3_PLF_138_net_1, \b7_vFW_PlM[252] , 
        \b7_vFW_PlM[12] , b3_PLF_137_net_1, \b7_vFW_PlM[141] , 
        \b7_vFW_PlM[30] , b3_PLF_136_net_1, \b7_vFW_PlM[286] , 
        \b7_vFW_PlM[175] , b3_PLF_135_net_1, \b7_vFW_PlM[304] , 
        \b7_vFW_PlM[48] , b3_PLF_134_net_1, \b7_vFW_PlM[177] , 
        \b7_vFW_PlM[50] , b3_PLF_133_net_1, \b7_vFW_PlM[306] , 
        \b7_vFW_PlM[179] , b3_PLF_132_net_1, \b7_vFW_PlM[308] , 
        \b7_vFW_PlM[52] , b3_PLF_131_net_1, \b7_vFW_PlM[181] , 
        \b7_vFW_PlM[54] , b3_PLF_130_net_1, \b7_vFW_PlM[310] , 
        \b7_vFW_PlM[183] , b3_PLF_129_net_1, \b7_vFW_PlM[312] , 
        \b7_vFW_PlM[56] , b3_PLF_128_net_1, \b7_vFW_PlM[185] , 
        \b7_vFW_PlM[74] , b3_PLF_127_net_1, \b7_vFW_PlM[347] , 
        \b7_vFW_PlM[91] , b3_PLF_126_net_1, \b7_vFW_PlM[236] , 
        \b7_vFW_PlM[125] , b3_PLF_125_net_1, \b7_vFW_PlM[365] , 
        \b7_vFW_PlM[270] , b3_PLF_124_net_1, \b7_vFW_PlM[159] , 
        \b7_vFW_PlM[32] , b3_PLF_123_net_1, \b7_vFW_PlM[288] , 
        \b7_vFW_PlM[161] , b3_PLF_122_net_1, \b7_vFW_PlM[290] , 
        \b7_vFW_PlM[34] , b3_PLF_121_net_1, \b7_vFW_PlM[163] , 
        \b7_vFW_PlM[36] , b3_PLF_120_net_1, \b7_vFW_PlM[292] , 
        \b7_vFW_PlM[165] , b3_PLF_119_net_1, \b7_vFW_PlM[294] , 
        \b7_vFW_PlM[38] , b3_PLF_118_net_1, \b7_vFW_PlM[167] , 
        \b7_vFW_PlM[40] , b3_PLF_117_net_1, \b7_vFW_PlM[296] , 
        \b7_vFW_PlM[169] , b3_PLF_116_net_1, \b7_vFW_PlM[75] , 
        \b7_vFW_PlM[58] , b3_PLF_115_net_1, \b7_vFW_PlM[331] , 
        \b7_vFW_PlM[220] , b3_PLF_114_net_1, \b7_vFW_PlM[109] , 
        \b7_vFW_PlM[14] , b3_PLF_113_net_1, \b7_vFW_PlM[254] , 
        \b7_vFW_PlM[143] , b3_PLF_112_net_1, \b7_vFW_PlM[272] , 
        \b7_vFW_PlM[16] , b3_PLF_111_net_1, \b7_vFW_PlM[145] , 
        \b7_vFW_PlM[18] , b3_PLF_110_net_1, \b7_vFW_PlM[274] , 
        \b7_vFW_PlM[147] , b3_PLF_109_net_1, \b7_vFW_PlM[276] , 
        \b7_vFW_PlM[20] , b3_PLF_108_net_1, \b7_vFW_PlM[149] , 
        \b7_vFW_PlM[22] , b3_PLF_107_net_1, \b7_vFW_PlM[278] , 
        \b7_vFW_PlM[151] , b3_PLF_106_net_1, \b7_vFW_PlM[280] , 
        \b7_vFW_PlM[24] , b3_PLF_105_net_1, \b7_vFW_PlM[153] , 
        \b7_vFW_PlM[42] , b3_PLF_104_net_1, \b7_vFW_PlM[315] , 
        \b7_vFW_PlM[59] , b3_PLF_103_net_1, \b7_vFW_PlM[204] , 
        \b7_vFW_PlM[93] , b3_PLF_102_net_1, \b7_vFW_PlM[349] , 
        \b7_vFW_PlM[238] , b3_PLF_101_net_1, \b7_vFW_PlM[127] , 
        \b7_vFW_PlM[0] , b3_PLF_100_net_1, \b7_vFW_PlM[256] , 
        \b7_vFW_PlM[129] , b3_PLF_99_net_1, \b7_vFW_PlM[258] , 
        \b7_vFW_PlM[2] , b3_PLF_98_net_1, \b7_vFW_PlM[131] , 
        \b7_vFW_PlM[4] , b3_PLF_97_net_1, \b7_vFW_PlM[260] , 
        \b7_vFW_PlM[133] , b3_PLF_96_net_1, \b7_vFW_PlM[262] , 
        \b7_vFW_PlM[6] , b3_PLF_95_net_1, \b7_vFW_PlM[135] , 
        \b7_vFW_PlM[8] , b3_PLF_94_net_1, \b7_vFW_PlM[264] , 
        \b7_vFW_PlM[137] , b3_PLF_93_net_1, \b7_vFW_PlM[43] , 
        \b7_vFW_PlM[26] , b3_PLF_92_net_1, \b7_vFW_PlM[299] , 
        \b7_vFW_PlM[188] , b3_PLF_91_net_1, \b7_vFW_PlM[333] , 
        \b7_vFW_PlM[77] , b3_PLF_90_net_1, \b7_vFW_PlM[222] , 
        \b7_vFW_PlM[111] , b3_PLF_89_net_1, \b7_vFW_PlM[367] , 
        \b7_vFW_PlM[240] , b3_PLF_88_net_1, \b7_vFW_PlM[369] , 
        \b7_vFW_PlM[113] , b3_PLF_87_net_1, \b7_vFW_PlM[242] , 
        \b7_vFW_PlM[115] , b3_PLF_86_net_1, \b7_vFW_PlM[371] , 
        \b7_vFW_PlM[244] , b3_PLF_85_net_1, \b7_vFW_PlM[373] , 
        \b7_vFW_PlM[117] , b3_PLF_84_net_1, \b7_vFW_PlM[246] , 
        \b7_vFW_PlM[119] , b3_PLF_83_net_1, \b7_vFW_PlM[375] , 
        \b7_vFW_PlM[248] , b3_PLF_82_net_1, \b7_vFW_PlM[361] , 
        \b7_vFW_PlM[121] , b3_PLF_81_net_1, \b7_vFW_PlM[266] , 
        \b7_vFW_PlM[27] , b3_PLF_80_net_1, \b7_vFW_PlM[283] , 
        \b7_vFW_PlM[172] , b3_PLF_79_net_1, \b7_vFW_PlM[317] , 
        \b7_vFW_PlM[61] , b3_PLF_78_net_1, \b7_vFW_PlM[206] , 
        \b7_vFW_PlM[95] , b3_PLF_77_net_1, \b7_vFW_PlM[351] , 
        \b7_vFW_PlM[224] , b3_PLF_76_net_1, \b7_vFW_PlM[353] , 
        \b7_vFW_PlM[97] , b3_PLF_75_net_1, \b7_vFW_PlM[226] , 
        \b7_vFW_PlM[99] , b3_PLF_74_net_1, \b7_vFW_PlM[355] , 
        \b7_vFW_PlM[228] , b3_PLF_73_net_1, \b7_vFW_PlM[357] , 
        \b7_vFW_PlM[101] , b3_PLF_72_net_1, \b7_vFW_PlM[230] , 
        \b7_vFW_PlM[103] , b3_PLF_71_net_1, \b7_vFW_PlM[359] , 
        \b7_vFW_PlM[232] , b3_PLF_70_net_1, \b7_vFW_PlM[105] , 
        \b7_vFW_PlM[10] , b3_PLF_69_net_1, \b7_vFW_PlM[250] , 
        \b7_vFW_PlM[11] , b3_PLF_68_net_1, \b7_vFW_PlM[267] , 
        \b7_vFW_PlM[156] , b3_PLF_67_net_1, \b7_vFW_PlM[301] , 
        \b7_vFW_PlM[45] , b3_PLF_66_net_1, \b7_vFW_PlM[190] , 
        \b7_vFW_PlM[79] , b3_PLF_65_net_1, \b7_vFW_PlM[335] , 
        \b7_vFW_PlM[208] , b3_PLF_64_net_1, \b7_vFW_PlM[337] , 
        \b7_vFW_PlM[81] , b3_PLF_63_net_1, \b7_vFW_PlM[210] , 
        \b7_vFW_PlM[83] , b3_PLF_62_net_1, \b7_vFW_PlM[339] , 
        \b7_vFW_PlM[212] , b3_PLF_61_net_1, \b7_vFW_PlM[341] , 
        \b7_vFW_PlM[85] , b3_PLF_60_net_1, \b7_vFW_PlM[214] , 
        \b7_vFW_PlM[87] , b3_PLF_59_net_1, \b7_vFW_PlM[343] , 
        \b7_vFW_PlM[216] , b3_PLF_58_net_1, \b7_vFW_PlM[345] , 
        \b7_vFW_PlM[89] , b3_PLF_57_net_1, \b7_vFW_PlM[362] , 
        \b7_vFW_PlM[234] , b3_PLF_56_net_1, \b7_vFW_PlM[251] , 
        \b7_vFW_PlM[140] , b3_PLF_55_net_1, \b7_vFW_PlM[285] , 
        \b7_vFW_PlM[29] , b3_PLF_54_net_1, \b7_vFW_PlM[174] , 
        \b7_vFW_PlM[63] , b3_PLF_53_net_1, \b7_vFW_PlM[319] , 
        \b7_vFW_PlM[192] , b3_PLF_52_net_1, \b7_vFW_PlM[321] , 
        \b7_vFW_PlM[65] , b3_PLF_51_net_1, \b7_vFW_PlM[194] , 
        \b7_vFW_PlM[67] , b3_PLF_50_net_1, \b7_vFW_PlM[323] , 
        \b7_vFW_PlM[196] , b3_PLF_49_net_1, \b7_vFW_PlM[325] , 
        \b7_vFW_PlM[69] , b3_PLF_48_net_1, \b7_vFW_PlM[198] , 
        \b7_vFW_PlM[71] , b3_PLF_47_net_1, \b7_vFW_PlM[327] , 
        \b7_vFW_PlM[200] , b3_PLF_46_net_1, \b7_vFW_PlM[329] , 
        \b7_vFW_PlM[73] , b3_PLF_45_net_1, \b7_vFW_PlM[346] , 
        \b7_vFW_PlM[218] , b3_PLF_44_net_1, \b7_vFW_PlM[235] , 
        \b7_vFW_PlM[124] , b3_PLF_43_net_1, \b7_vFW_PlM[269] , 
        \b7_vFW_PlM[13] , b3_PLF_42_net_1, \b7_vFW_PlM[158] , 
        \b7_vFW_PlM[47] , b3_PLF_41_net_1, \b7_vFW_PlM[303] , 
        \b7_vFW_PlM[176] , b3_PLF_40_net_1, \b7_vFW_PlM[305] , 
        \b7_vFW_PlM[49] , b3_PLF_39_net_1, \b7_vFW_PlM[178] , 
        \b7_vFW_PlM[51] , b3_PLF_38_net_1, \b7_vFW_PlM[307] , 
        \b7_vFW_PlM[180] , b3_PLF_37_net_1, \b7_vFW_PlM[309] , 
        \b7_vFW_PlM[53] , b3_PLF_36_net_1, \b7_vFW_PlM[182] , 
        \b7_vFW_PlM[55] , b3_PLF_35_net_1, \b7_vFW_PlM[311] , 
        \b7_vFW_PlM[184] , b3_PLF_34_net_1, \b7_vFW_PlM[313] , 
        \b7_vFW_PlM[57] , b3_PLF_33_net_1, \b7_vFW_PlM[330] , 
        \b7_vFW_PlM[202] , b3_PLF_32_net_1, \b7_vFW_PlM[219] , 
        \b7_vFW_PlM[108] , b3_PLF_31_net_1, \b7_vFW_PlM[364] , 
        \b7_vFW_PlM[253] , b3_PLF_30_net_1, \b7_vFW_PlM[142] , 
        \b7_vFW_PlM[31] , b3_PLF_29_net_1, \b7_vFW_PlM[287] , 
        \b7_vFW_PlM[160] , b3_PLF_28_net_1, \b7_vFW_PlM[289] , 
        \b7_vFW_PlM[33] , b3_PLF_27_net_1, \b7_vFW_PlM[162] , 
        \b7_vFW_PlM[35] , b3_PLF_26_net_1, \b7_vFW_PlM[291] , 
        \b7_vFW_PlM[164] , b3_PLF_25_net_1, \b7_vFW_PlM[293] , 
        \b7_vFW_PlM[37] , b3_PLF_24_net_1, \b7_vFW_PlM[166] , 
        \b7_vFW_PlM[39] , b3_PLF_23_net_1, \b7_vFW_PlM[295] , 
        \b7_vFW_PlM[168] , b3_PLF_22_net_1, \b7_vFW_PlM[297] , 
        \b7_vFW_PlM[41] , b3_PLF_21_net_1, \b7_vFW_PlM[314] , 
        \b7_vFW_PlM[186] , b3_PLF_20_net_1, \b7_vFW_PlM[203] , 
        \b7_vFW_PlM[92] , b3_PLF_19_net_1, \b7_vFW_PlM[348] , 
        \b7_vFW_PlM[237] , b3_PLF_18_net_1, \b7_vFW_PlM[126] , 
        \b7_vFW_PlM[15] , b3_PLF_17_net_1, \b7_vFW_PlM[271] , 
        \b7_vFW_PlM[144] , b3_PLF_16_net_1, \b7_vFW_PlM[273] , 
        \b7_vFW_PlM[17] , b3_PLF_15_net_1, \b7_vFW_PlM[146] , 
        \b7_vFW_PlM[19] , b3_PLF_14_net_1, \b7_vFW_PlM[275] , 
        \b7_vFW_PlM[148] , b3_PLF_13_net_1, \b7_vFW_PlM[277] , 
        \b7_vFW_PlM[21] , b3_PLF_12_net_1, \b7_vFW_PlM[150] , 
        \b7_vFW_PlM[23] , b3_PLF_11_net_1, \b7_vFW_PlM[279] , 
        \b7_vFW_PlM[152] , b3_PLF_10_net_1, \b7_vFW_PlM[281] , 
        \b7_vFW_PlM[25] , b3_PLF_9_net_1, \b7_vFW_PlM[298] , 
        \b7_vFW_PlM[170] , b3_PLF_8_net_1, \b7_vFW_PlM[187] , 
        \b7_vFW_PlM[76] , b3_PLF_7_net_1, \b7_vFW_PlM[332] , 
        \b7_vFW_PlM[221] , b3_PLF_6_net_1, \b7_vFW_PlM[366] , 
        \b7_vFW_PlM[110] , b3_PLF_5_net_1, \b7_vFW_PlM[255] , 
        \b7_vFW_PlM[128] , b3_PLF_4_net_1, \b7_vFW_PlM[130] , 
        \b7_vFW_PlM[3] , b3_PLF_2_net_1, \b7_vFW_PlM[259] , 
        \b7_vFW_PlM[132] , b3_PLF_1_net_1, \b7_vFW_PlM[261] , 
        \b7_vFW_PlM[5] , b3_PLF_0_net_1, b8_jAA_KlCO_0_sqmuxa_6_net_1, 
        m9_e_6, m9_e_5, \b7_vFW_PlM[154] , b3_PLF_281_net_1, 
        \b7_vFW_PlM[257] , b3_PLF_190_net_1, \b7_vFW_PlM[134] , 
        b3_PLF_188_net_1, b8_jAA_KlCO_0_sqmuxa_8_net_1, 
        un1_b13_PLF_2grFt_FH911_i_a2_0_2, b3_PLF_328_net_1, 
        b3_PLF_327_net_1, b3_PLF_326_net_1, b3_PLF_325_net_1, 
        b3_PLF_324_net_1, b3_PLF_323_net_1, b3_PLF_322_net_1, 
        b3_PLF_321_net_1, b3_PLF_320_net_1, b3_PLF_319_net_1, 
        b3_PLF_318_net_1, b3_PLF_317_net_1, b3_PLF_316_net_1, 
        b3_PLF_315_net_1, b3_PLF_314_net_1, b3_PLF_313_net_1, 
        b3_PLF_312_net_1, b3_PLF_311_net_1, b3_PLF_310_net_1, 
        b3_PLF_309_net_1, b3_PLF_308_net_1, b3_PLF_307_net_1, 
        b3_PLF_306_net_1, b3_PLF_305_net_1, b3_PLF_304_net_1, 
        b3_PLF_303_net_1, b3_PLF_302_net_1, b3_PLF_301_net_1, 
        b3_PLF_300_net_1, b3_PLF_299_net_1, b3_PLF_298_net_1, 
        b3_PLF_297_net_1, b3_PLF_296_net_1, b3_PLF_295_net_1, 
        b3_PLF_294_net_1, b3_PLF_293_net_1, b3_PLF_292_net_1, 
        b3_PLF_291_net_1, b3_PLF_290_net_1, b3_PLF_289_net_1, 
        b3_PLF_288_net_1, b3_PLF_287_net_1, b3_PLF_286_net_1, 
        b3_PLF_285_net_1, b3_PLF_284_net_1, b3_PLF_330_net_1, 
        b3_PLF_364_net_1, b3_PLF_363_net_1, b3_PLF_362_net_1, 
        b3_PLF_361_net_1, b3_PLF_360_net_1, b3_PLF_359_net_1, 
        b3_PLF_358_net_1, b3_PLF_357_net_1, b3_PLF_356_net_1, 
        b3_PLF_355_net_1, b3_PLF_354_net_1, b3_PLF_353_net_1, 
        b3_PLF_373_net_1, b3_PLF_372_net_1, b3_PLF_371_net_1, N_21, 
        un1_b5_OvyH3;
    
    SLE \genblk9.b7_nYJ_BFM[210]  (.D(\b7_nYJ_BFM[209] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[210] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_94 (.A(\b7_nYJ_BFM[136] ), .B(
        \b7_nYJ_BFM[9] ), .C(\b7_vFW_PlM[135] ), .D(\b7_vFW_PlM[8] ), 
        .Y(b3_PLF_94_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_108 (.A(\b7_nYJ_BFM[277] ), .B(
        \b7_nYJ_BFM[21] ), .C(\b7_vFW_PlM[276] ), .D(\b7_vFW_PlM[20] ), 
        .Y(b3_PLF_108_net_1));
    SLE \genblk9.b7_nYJ_BFM[34]  (.D(\b7_nYJ_BFM[33] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[34] ));
    SLE \genblk9.b7_nYJ_BFM[202]  (.D(\b7_nYJ_BFM[201] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[202] ));
    SLE \genblk9.b7_nYJ_BFM[314]  (.D(\b7_nYJ_BFM[313] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[314] ));
    SLE \genblk9.b7_nYJ_BFM[48]  (.D(\b7_nYJ_BFM[47] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[48] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_70 (.A(\b7_nYJ_BFM[360] ), .B(
        \b7_nYJ_BFM[233] ), .C(\b7_vFW_PlM[359] ), .D(
        \b7_vFW_PlM[232] ), .Y(b3_PLF_70_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_27 (.A(\b7_nYJ_BFM[290] ), .B(
        \b7_nYJ_BFM[34] ), .C(\b7_vFW_PlM[289] ), .D(\b7_vFW_PlM[33] ), 
        .Y(b3_PLF_27_net_1));
    SLE \genblk9.b7_nYJ_BFM[158]  (.D(\b7_nYJ_BFM[157] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[158] ));
    SLE \genblk9.b7_nYJ_BFM[27]  (.D(\b7_nYJ_BFM[26] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[27] ));
    SLE \genblk9.b9_v_mzCDYXs[3]  (.D(b9_v_mzCDYXs), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[3] ));
    SLE \genblk9.b7_nYJ_BFM[95]  (.D(\b7_nYJ_BFM[94] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[95] ));
    SLE \genblk9.b7_nYJ_BFM[294]  (.D(\b7_nYJ_BFM[293] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[294] ));
    SLE \genblk9.b7_nYJ_BFM[167]  (.D(\b7_nYJ_BFM[166] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[167] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_138 (.A(\b7_nYJ_BFM[108] ), .B(
        \b7_nYJ_BFM[91] ), .C(\b7_vFW_PlM[107] ), .D(\b7_vFW_PlM[90] ), 
        .Y(b3_PLF_138_net_1));
    SLE \genblk9.b7_nYJ_BFM[147]  (.D(\b7_nYJ_BFM[146] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[147] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[0]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_0_S), .Y(b12_2_St6KCa_jHv));
    SLE \genblk9.b7_nYJ_BFM[71]  (.D(\b7_nYJ_BFM[70] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[71] ));
    SLE \genblk9.b7_nYJ_BFM[322]  (.D(\b7_nYJ_BFM[321] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[322] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[6]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_6_S), .Y(b12_2_St6KCa_jHv_5));
    SLE \genblk9.b7_nYJ_BFM[280]  (.D(\b7_nYJ_BFM[279] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[280] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_8 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[8]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_7_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_8_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_8_net_1));
    SLE \genblk9.b7_nYJ_BFM[321]  (.D(\b7_nYJ_BFM[320] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[321] ));
    SLE \genblk9.b7_nYJ_BFM[298]  (.D(\b7_nYJ_BFM[297] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[298] ));
    SLE \genblk9.b7_nYJ_BFM[227]  (.D(\b7_nYJ_BFM[226] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[227] ));
    SLE \genblk9.b7_nYJ_BFM[61]  (.D(\b7_nYJ_BFM[60] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[61] ));
    SLE \genblk9.b7_nYJ_BFM[367]  (.D(\b7_nYJ_BFM[366] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[367] ));
    SLE \genblk9.b7_nYJ_BFM[347]  (.D(\b7_nYJ_BFM[346] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[347] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNI4UHH6[5]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[5] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_4), .S(\b9_v_mzCDYXs_RNI4UHH6_S[5] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_5));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_73 (.A(\b7_nYJ_BFM[356] ), .B(
        \b7_nYJ_BFM[229] ), .C(\b7_vFW_PlM[355] ), .D(
        \b7_vFW_PlM[228] ), .Y(b3_PLF_73_net_1));
    SLE \genblk9.b7_nYJ_BFM[336]  (.D(\b7_nYJ_BFM[335] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[336] ));
    SLE \genblk9.b7_nYJ_BFM[372]  (.D(\b7_nYJ_BFM[371] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[372] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_117 (.A(\b7_nYJ_BFM[168] ), .B(
        \b7_nYJ_BFM[41] ), .C(\b7_vFW_PlM[167] ), .D(\b7_vFW_PlM[40] ), 
        .Y(b3_PLF_117_net_1));
    CFG2 #( .INIT(4'h8) )  \genblk9.un1_b4_BVmQ[265]  (.A(
        \b7_vFW_PlM[265] ), .B(\b7_nYJ_BFM[266] ), .Y(
        \un1_b4_BVmQ[265] ));
    SLE \genblk9.b7_nYJ_BFM[368]  (.D(\b7_nYJ_BFM[367] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[368] ));
    SLE \genblk9.b7_nYJ_BFM[201]  (.D(\b7_nYJ_BFM[200] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[201] ));
    SLE \genblk9.b7_nYJ_BFM[348]  (.D(\b7_nYJ_BFM[347] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[348] ));
    SLE \genblk9.b7_nYJ_BFM[371]  (.D(\b7_nYJ_BFM[370] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[371] ));
    SLE \genblk9.b7_nYJ_BFM[199]  (.D(\b7_nYJ_BFM[198] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[199] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNILNNS6[6]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[6] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_5), .S(\b9_v_mzCDYXs_RNILNNS6_S[6] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_6));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_24 (.A(\b7_nYJ_BFM[294] ), .B(
        \b7_nYJ_BFM[38] ), .C(\b7_vFW_PlM[293] ), .D(\b7_vFW_PlM[37] ), 
        .Y(b3_PLF_24_net_1));
    SLE \genblk9.b7_nYJ_BFM[277]  (.D(\b7_nYJ_BFM[276] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[277] ));
    SLE \genblk9.b7_nYJ_BFM[230]  (.D(\b7_nYJ_BFM[229] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[230] ));
    SLE \genblk9.b9_v_mzCDYXs[2]  (.D(b9_v_mzCDYXs_0), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[2] ));
    SLE \genblk9.b7_nYJ_BFM[80]  (.D(\b7_nYJ_BFM[79] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[80] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_15 (.A(\b7_nYJ_BFM[274] ), .B(
        \b7_nYJ_BFM[18] ), .C(\b7_vFW_PlM[273] ), .D(\b7_vFW_PlM[17] ), 
        .Y(b3_PLF_15_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_300 (.A(b3_PLF_72_net_1), .B(
        b3_PLF_71_net_1), .C(b3_PLF_70_net_1), .D(b3_PLF_69_net_1), .Y(
        b3_PLF_300_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_328 (.A(b3_PLF_184_net_1), .B(
        b3_PLF_183_net_1), .C(b3_PLF_182_net_1), .D(b3_PLF_181_net_1), 
        .Y(b3_PLF_328_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_31 (.A(\b7_nYJ_BFM[220] ), .B(
        \b7_nYJ_BFM[109] ), .C(\b7_vFW_PlM[219] ), .D(
        \b7_vFW_PlM[108] ), .Y(b3_PLF_31_net_1));
    SLE \genblk9.b7_nYJ_BFM[312]  (.D(\b7_nYJ_BFM[311] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[312] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_112 (.A(\b7_nYJ_BFM[255] ), .B(
        \b7_nYJ_BFM[144] ), .C(\b7_vFW_PlM[254] ), .D(
        \b7_vFW_PlM[143] ), .Y(b3_PLF_112_net_1));
    SLE \genblk9.b7_nYJ_BFM[120]  (.D(\b7_nYJ_BFM[119] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[120] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_18 (.A(\b7_nYJ_BFM[349] ), .B(
        \b7_nYJ_BFM[238] ), .C(\b7_vFW_PlM[348] ), .D(
        \b7_vFW_PlM[237] ), .Y(b3_PLF_18_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_55 (.A(\b7_nYJ_BFM[252] ), .B(
        \b7_nYJ_BFM[141] ), .C(\b7_vFW_PlM[251] ), .D(
        \b7_vFW_PlM[140] ), .Y(b3_PLF_55_net_1));
    SLE \genblk9.b7_nYJ_BFM[334]  (.D(\b7_nYJ_BFM[333] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[334] ));
    SLE \b12_PSyi_KyDbLbb[7]  (.D(\b12_2_St6KCa_jHv[7]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[7]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[91]  (.D(\b7_nYJ_BFM[90] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[91] ));
    SLE \genblk9.b7_nYJ_BFM[311]  (.D(\b7_nYJ_BFM[310] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[311] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_42 (.A(\b7_nYJ_BFM[270] ), .B(
        \b7_nYJ_BFM[14] ), .C(\b7_vFW_PlM[269] ), .D(\b7_vFW_PlM[13] ), 
        .Y(b3_PLF_42_net_1));
    SLE \genblk9.b7_nYJ_BFM[217]  (.D(\b7_nYJ_BFM[216] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[217] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_58 (.A(\b7_nYJ_BFM[344] ), .B(
        \b7_nYJ_BFM[217] ), .C(\b7_vFW_PlM[343] ), .D(
        \b7_vFW_PlM[216] ), .Y(b3_PLF_58_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_324 (.A(b3_PLF_168_net_1), .B(
        b3_PLF_167_net_1), .C(b3_PLF_166_net_1), .D(b3_PLF_165_net_1), 
        .Y(b3_PLF_324_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_303 (.A(b3_PLF_84_net_1), .B(
        b3_PLF_83_net_1), .C(b3_PLF_82_net_1), .D(b3_PLF_81_net_1), .Y(
        b3_PLF_303_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[8]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNIQD3J7_S[8] ), .Y(b9_v_mzCDYXs_4));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b7_nYJ_BFM_RNI95U74[383]  (.A(
        b8_nYJ_TqLY), .B(N_24_mux), .C(IICE_comm2iice_10), .D(
        b10_OFWNT9khFt), .Y(\b7_nYJ_BFM_RNI95U74[383] ));
    SLE \genblk9.b7_nYJ_BFM[195]  (.D(\b7_nYJ_BFM[194] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[195] ));
    SLE \genblk9.b7_nYJ_BFM[170]  (.D(\b7_nYJ_BFM[169] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[170] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_4 (.A(\b7_nYJ_BFM[256] ), .B(
        \b7_nYJ_BFM[129] ), .C(\b7_vFW_PlM[255] ), .D(
        \b7_vFW_PlM[128] ), .Y(b3_PLF_4_net_1));
    SLE \genblk9.b7_nYJ_BFM[369]  (.D(\b7_nYJ_BFM[368] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[369] ));
    SLE \genblk9.b7_nYJ_BFM[349]  (.D(\b7_nYJ_BFM[348] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[349] ));
    SLE \genblk9.b7_nYJ_BFM[303]  (.D(\b7_nYJ_BFM[302] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[303] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_177 (.A(\b7_nYJ_BFM[373] ), .B(
        \b7_nYJ_BFM[117] ), .C(\b7_vFW_PlM[372] ), .D(
        \b7_vFW_PlM[116] ), .Y(b3_PLF_177_net_1));
    SLE \genblk9.b7_nYJ_BFM[56]  (.D(\b7_nYJ_BFM[55] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[56] ));
    SLE \genblk9.b7_nYJ_BFM[252]  (.D(\b7_nYJ_BFM[251] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[252] ));
    SLE \genblk9.b7_nYJ_BFM[193]  (.D(\b7_nYJ_BFM[192] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[193] ));
    SLE \genblk9.b7_nYJ_BFM[12]  (.D(\b7_nYJ_BFM[11] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[12] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_330 (.A(b3_PLF_1_net_1), .B(
        b3_PLF_2_net_1), .C(b3_PLF_284_net_1), .D(b3_PLF_190_net_1), 
        .Y(b3_PLF_330_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_361 (.A(b3_PLF_316_net_1), .B(
        b3_PLF_315_net_1), .C(b3_PLF_314_net_1), .D(b3_PLF_313_net_1), 
        .Y(b3_PLF_361_net_1));
    SLE \genblk9.b7_nYJ_BFM[265]  (.D(\b7_nYJ_BFM[264] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[265] ));
    SLE \genblk9.b7_nYJ_BFM[245]  (.D(\b7_nYJ_BFM[244] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[245] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_322 (.A(b3_PLF_160_net_1), .B(
        b3_PLF_159_net_1), .C(b3_PLF_158_net_1), .D(b3_PLF_157_net_1), 
        .Y(b3_PLF_322_net_1));
    SLE \genblk9.b7_nYJ_BFM[36]  (.D(\b7_nYJ_BFM[35] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[36] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_166 (.A(\b7_nYJ_BFM[228] ), .B(
        \b7_nYJ_BFM[101] ), .C(\b7_vFW_PlM[227] ), .D(
        \b7_vFW_PlM[100] ), .Y(b3_PLF_166_net_1));
    SLE \genblk9.b7_nYJ_BFM[382]  (.D(\b7_nYJ_BFM[381] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[382] ));
    SLE \genblk9.b7_nYJ_BFM[110]  (.D(\b7_nYJ_BFM[109] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[110] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_37 (.A(\b7_nYJ_BFM[308] ), .B(
        \b7_nYJ_BFM[181] ), .C(\b7_vFW_PlM[307] ), .D(
        \b7_vFW_PlM[180] ), .Y(b3_PLF_37_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_172 (.A(\b7_nYJ_BFM[156] ), .B(
        \b7_nYJ_BFM[45] ), .C(\b7_vFW_PlM[155] ), .D(\b7_vFW_PlM[44] ), 
        .Y(b3_PLF_172_net_1));
    SLE \genblk9.b7_nYJ_BFM[194]  (.D(\b7_nYJ_BFM[193] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[194] ));
    SLE \genblk9.b7_nYJ_BFM[381]  (.D(\b7_nYJ_BFM[380] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[381] ));
    SLE \genblk9.b7_nYJ_BFM[287]  (.D(\b7_nYJ_BFM[286] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[287] ));
    SLE \genblk9.b7_nYJ_BFM[206]  (.D(\b7_nYJ_BFM[205] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[206] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_128 (.A(\b7_nYJ_BFM[313] ), .B(
        \b7_nYJ_BFM[57] ), .C(\b7_vFW_PlM[312] ), .D(\b7_vFW_PlM[56] ), 
        .Y(b3_PLF_128_net_1));
    SLE \genblk9.b7_nYJ_BFM[161]  (.D(\b7_nYJ_BFM[160] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[161] ));
    SLE \b12_2_St6KCa_jHv[5]  (.D(b12_2_St6KCa_jHv_4), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[5]_net_1 ));
    SLE \genblk9.b9_v_mzCDYXs[4]  (.D(b9_v_mzCDYXs_8), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[4] ));
    SLE \genblk9.b7_nYJ_BFM[141]  (.D(\b7_nYJ_BFM[140] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[141] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[3]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_3_S), .Y(b12_2_St6KCa_jHv_2));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_147 (.A(\b7_nYJ_BFM[303] ), .B(
        \b7_nYJ_BFM[47] ), .C(\b7_vFW_PlM[302] ), .D(\b7_vFW_PlM[46] ), 
        .Y(b3_PLF_147_net_1));
    SLE \genblk9.b7_nYJ_BFM[332]  (.D(\b7_nYJ_BFM[331] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[332] ));
    SLE \b8_FZFFLXYE[4]  (.D(\b12_2_St6KCa_jHv[4]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[4]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[331]  (.D(\b7_nYJ_BFM[330] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[331] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_72 (.A(\b7_nYJ_BFM[358] ), .B(
        \b7_nYJ_BFM[102] ), .C(\b7_vFW_PlM[357] ), .D(
        \b7_vFW_PlM[101] ), .Y(b3_PLF_72_net_1));
    SLE \b8_FZFFLXYE[0]  (.D(\b12_2_St6KCa_jHv[0]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[0]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[237]  (.D(\b7_nYJ_BFM[236] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[237] ));
    SLE \genblk9.b9_v_mzCDYXs[7]  (.D(b9_v_mzCDYXs_5), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[7] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_165 (.A(\b7_nYJ_BFM[357] ), .B(
        \b7_nYJ_BFM[230] ), .C(\b7_vFW_PlM[356] ), .D(
        \b7_vFW_PlM[229] ), .Y(b3_PLF_165_net_1));
    SLE \genblk9.b7_nYJ_BFM[224]  (.D(\b7_nYJ_BFM[223] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[224] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[7]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNI7IT77_S[7] ), .Y(b9_v_mzCDYXs_5));
    SLE \genblk9.b7_nYJ_BFM[251]  (.D(\b7_nYJ_BFM[250] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[251] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_34 (.A(\b7_nYJ_BFM[312] ), .B(
        \b7_nYJ_BFM[185] ), .C(\b7_vFW_PlM[311] ), .D(
        \b7_vFW_PlM[184] ), .Y(b3_PLF_34_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_142 (.A(\b7_nYJ_BFM[325] ), .B(
        \b7_nYJ_BFM[198] ), .C(\b7_vFW_PlM[324] ), .D(
        \b7_vFW_PlM[197] ), .Y(b3_PLF_142_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_7 (.A(\b7_nYJ_BFM[188] ), .B(
        \b7_nYJ_BFM[77] ), .C(\b7_vFW_PlM[187] ), .D(\b7_vFW_PlM[76] ), 
        .Y(b3_PLF_7_net_1));
    SLE \genblk9.b7_nYJ_BFM[180]  (.D(\b7_nYJ_BFM[179] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[180] ));
    SLE \genblk9.b7_nYJ_BFM[293]  (.D(\b7_nYJ_BFM[292] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[293] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_99 (.A(\b7_nYJ_BFM[257] ), .B(
        \b7_nYJ_BFM[130] ), .C(\b7_vFW_PlM[256] ), .D(
        \b7_vFW_PlM[129] ), .Y(b3_PLF_99_net_1));
    SLE \b8_FZFFLXYE[2]  (.D(\b12_2_St6KCa_jHv[2]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[2]_net_1 ));
    SLE \b8_FZFFLXYE[8]  (.D(\b12_2_St6KCa_jHv[8]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[8]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[228]  (.D(\b7_nYJ_BFM[227] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[228] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_307 (.A(b3_PLF_100_net_1), .B(
        b3_PLF_99_net_1), .C(b3_PLF_98_net_1), .D(b3_PLF_97_net_1), .Y(
        b3_PLF_307_net_1));
    SLE \genblk9.b7_nYJ_BFM[274]  (.D(\b7_nYJ_BFM[273] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[274] ));
    SLE \genblk9.b7_nYJ_BFM[192]  (.D(\b7_nYJ_BFM[191] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[192] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_1 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[1]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_0_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_1_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_1_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_287 (.A(b3_PLF_20_net_1), .B(
        b3_PLF_19_net_1), .C(b3_PLF_18_net_1), .D(b3_PLF_17_net_1), .Y(
        b3_PLF_287_net_1));
    GND GND (.Y(GND_net_1));
    SLE \genblk9.b7_nYJ_BFM[25]  (.D(\b7_nYJ_BFM[24] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[25] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_100 (.A(\b7_nYJ_BFM[128] ), .B(
        \b7_nYJ_BFM[1] ), .C(\b7_vFW_PlM[127] ), .D(\b7_vFW_PlM[0] ), 
        .Y(b3_PLF_100_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_r_RNO[9]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[9] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_8), .S(\b9_v_mzCDYXs_r_RNO_S[9] ), .Y()
        , .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNI7IT77[7]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[7] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_6), .S(\b9_v_mzCDYXs_RNI7IT77_S[7] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_7));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNI5E6R5[3]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[3] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_2), .S(\b9_v_mzCDYXs_RNI5E6R5_S[3] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_3));
    SLE \genblk9.b7_nYJ_BFM[166]  (.D(\b7_nYJ_BFM[165] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[166] ));
    SLE \genblk9.b7_nYJ_BFM[146]  (.D(\b7_nYJ_BFM[145] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[146] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_103 (.A(\b7_nYJ_BFM[316] ), .B(
        \b7_nYJ_BFM[60] ), .C(\b7_vFW_PlM[315] ), .D(\b7_vFW_PlM[59] ), 
        .Y(b3_PLF_103_net_1));
    SLE \genblk9.b7_nYJ_BFM[129]  (.D(\b7_nYJ_BFM[128] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[129] ));
    SLE \genblk9.b7_nYJ_BFM[72]  (.D(\b7_nYJ_BFM[71] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[72] ));
    SLE \genblk9.b7_nYJ_BFM[278]  (.D(\b7_nYJ_BFM[277] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[278] ));
    SLE \genblk9.b7_nYJ_BFM[130]  (.D(\b7_nYJ_BFM[129] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[130] ));
    SLE \genblk9.b7_nYJ_BFM[83]  (.D(\b7_nYJ_BFM[82] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[83] ));
    SLE \genblk9.b7_nYJ_BFM[214]  (.D(\b7_nYJ_BFM[213] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[214] ));
    SLE \genblk9.b7_nYJ_BFM[353]  (.D(\b7_nYJ_BFM[352] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[353] ));
    SLE \genblk9.b7_nYJ_BFM[19]  (.D(\b7_nYJ_BFM[18] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[19] ));
    SLE \genblk9.b7_nYJ_BFM[62]  (.D(\b7_nYJ_BFM[61] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[62] ));
    SLE \genblk9.b7_nYJ_BFM[179]  (.D(\b7_nYJ_BFM[178] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[179] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_355 (.A(b3_PLF_292_net_1), .B(
        b3_PLF_291_net_1), .C(b3_PLF_290_net_1), .D(b3_PLF_289_net_1), 
        .Y(b3_PLF_355_net_1));
    SLE \b12_2_St6KCa_jHv[0]  (.D(b12_2_St6KCa_jHv), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[0]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[320]  (.D(\b7_nYJ_BFM[319] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[320] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_320 (.A(b3_PLF_152_net_1), .B(
        b3_PLF_151_net_1), .C(b3_PLF_150_net_1), .D(b3_PLF_149_net_1), 
        .Y(b3_PLF_320_net_1));
    SLE \b12_2_St6KCa_jHv[6]  (.D(b12_2_St6KCa_jHv_5), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_161 (.A(\b7_nYJ_BFM[140] ), .B(
        \b7_nYJ_BFM[123] ), .C(\b7_vFW_PlM[139] ), .D(
        \b7_vFW_PlM[122] ), .Y(b3_PLF_161_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_156 (.A(\b7_nYJ_BFM[210] ), .B(
        \b7_nYJ_BFM[83] ), .C(\b7_vFW_PlM[209] ), .D(\b7_vFW_PlM[82] ), 
        .Y(b3_PLF_156_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_130 (.A(\b7_nYJ_BFM[182] ), .B(
        \b7_nYJ_BFM[55] ), .C(\b7_vFW_PlM[181] ), .D(\b7_vFW_PlM[54] ), 
        .Y(b3_PLF_130_net_1));
    SLE \genblk9.b7_nYJ_BFM[218]  (.D(\b7_nYJ_BFM[217] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[218] ));
    CFG3 #( .INIT(8'hFE) )  b3_PLF (.A(b3_PLF_373_net_1), .B(
        b3_PLF_372_net_1), .C(b3_PLF_371_net_1), .Y(b9_OFWNT9Mxf));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_133 (.A(\b7_nYJ_BFM[178] ), .B(
        \b7_nYJ_BFM[51] ), .C(\b7_vFW_PlM[177] ), .D(\b7_vFW_PlM[50] ), 
        .Y(b3_PLF_133_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_186 (.A(\b7_nYJ_BFM[137] ), .B(
        \b7_nYJ_BFM[10] ), .C(\b7_vFW_PlM[136] ), .D(\b7_vFW_PlM[9] ), 
        .Y(b3_PLF_186_net_1));
    SLE b9_PSyil9s_2 (.D(b11_PSyil9s_FMZ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b9_PSyil9s_2_net_1));
    SLE \genblk9.b7_nYJ_BFM[370]  (.D(\b7_nYJ_BFM[369] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[370] ));
    SLE \genblk9.b7_nYJ_BFM[40]  (.D(\b7_nYJ_BFM[39] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[40] ));
    SLE \genblk9.b7_nYJ_BFM[57]  (.D(\b7_nYJ_BFM[56] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[57] ));
    SLE \genblk9.b7_nYJ_BFM[125]  (.D(\b7_nYJ_BFM[124] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[125] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_323 (.A(b3_PLF_164_net_1), .B(
        b3_PLF_163_net_1), .C(b3_PLF_162_net_1), .D(b3_PLF_161_net_1), 
        .Y(b3_PLF_323_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_29 (.A(\b7_nYJ_BFM[143] ), .B(
        \b7_nYJ_BFM[32] ), .C(\b7_vFW_PlM[142] ), .D(\b7_vFW_PlM[31] ), 
        .Y(b3_PLF_29_net_1));
    SLE \genblk9.b7_nYJ_BFM[119]  (.D(\b7_nYJ_BFM[118] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[119] ));
    SLE \genblk9.b7_nYJ_BFM[123]  (.D(\b7_nYJ_BFM[122] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[123] ));
    SLE \genblk9.b7_nYJ_BFM[256]  (.D(\b7_nYJ_BFM[255] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[256] ));
    SLE \genblk9.b7_nYJ_BFM[37]  (.D(\b7_nYJ_BFM[36] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[37] ));
    CFG2 #( .INIT(4'hE) )  \genblk9.b7_nYJ_BFM_or[7]  (.A(
        N_850_a2_1_net_1), .B(b8_SoWGfWYY), .Y(\b7_nYJ_BFM_or[7] ));
    SLE \genblk9.b7_nYJ_BFM[21]  (.D(\b7_nYJ_BFM[20] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[21] ));
    SLE \genblk9.b7_nYJ_BFM[84]  (.D(\b7_nYJ_BFM[83] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[84] ));
    SLE \genblk9.b7_nYJ_BFM[175]  (.D(\b7_nYJ_BFM[174] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[175] ));
    SLE \genblk9.b7_nYJ_BFM[92]  (.D(\b7_nYJ_BFM[91] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[92] ));
    SLE \genblk9.b7_nYJ_BFM[284]  (.D(\b7_nYJ_BFM[283] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[284] ));
    SLE \genblk9.b7_nYJ_BFM[18]  (.D(\b7_nYJ_BFM[17] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[18] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[8]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_8_S), .Y(b12_2_St6KCa_jHv_7));
    SLE \genblk9.b7_nYJ_BFM[198]  (.D(\b7_nYJ_BFM[197] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[198] ));
    SLE \genblk9.b7_nYJ_BFM[173]  (.D(\b7_nYJ_BFM[172] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[173] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_155 (.A(\b7_nYJ_BFM[339] ), .B(
        \b7_nYJ_BFM[212] ), .C(\b7_vFW_PlM[338] ), .D(
        \b7_vFW_PlM[211] ), .Y(b3_PLF_155_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_114 (.A(\b7_nYJ_BFM[332] ), .B(
        \b7_nYJ_BFM[221] ), .C(\b7_vFW_PlM[331] ), .D(
        \b7_vFW_PlM[220] ), .Y(b3_PLF_114_net_1));
    SLE \genblk9.b7_nYJ_BFM[310]  (.D(\b7_nYJ_BFM[309] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[310] ));
    SLE \genblk9.b9_v_mzCDYXs[1]  (.D(b9_v_mzCDYXs_1), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[1] ));
    SLE \genblk9.b7_nYJ_BFM[124]  (.D(\b7_nYJ_BFM[123] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[124] ));
    SLE \genblk9.b7_nYJ_BFM[288]  (.D(\b7_nYJ_BFM[287] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[288] ));
    SLE \genblk9.b7_nYJ_BFM[107]  (.D(\b7_nYJ_BFM[106] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[107] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_169 (.A(\b7_nYJ_BFM[224] ), .B(
        \b7_nYJ_BFM[97] ), .C(\b7_vFW_PlM[223] ), .D(\b7_vFW_PlM[96] ), 
        .Y(b3_PLF_169_net_1));
    SLE \genblk9.b7_nYJ_BFM[234]  (.D(\b7_nYJ_BFM[233] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[234] ));
    SLE \genblk9.b7_nYJ_BFM[115]  (.D(\b7_nYJ_BFM[114] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[115] ));
    SLE \genblk9.b7_nYJ_BFM[174]  (.D(\b7_nYJ_BFM[173] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[174] ));
    SLE \genblk9.b7_nYJ_BFM[189]  (.D(\b7_nYJ_BFM[188] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[189] ));
    SLE \genblk9.b7_nYJ_BFM[113]  (.D(\b7_nYJ_BFM[112] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[113] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[4]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNIK5C66_S[4] ), .Y(b9_v_mzCDYXs_8));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_81 (.A(\b7_nYJ_BFM[362] ), .B(
        \b7_nYJ_BFM[122] ), .C(\b7_vFW_PlM[361] ), .D(
        \b7_vFW_PlM[121] ), .Y(b3_PLF_81_net_1));
    SLE \genblk9.b7_nYJ_BFM[307]  (.D(\b7_nYJ_BFM[306] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[307] ));
    SLE \genblk9.b7_nYJ_BFM[238]  (.D(\b7_nYJ_BFM[237] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[238] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_61 (.A(\b7_nYJ_BFM[340] ), .B(
        \b7_nYJ_BFM[213] ), .C(\b7_vFW_PlM[339] ), .D(
        \b7_vFW_PlM[212] ), .Y(b3_PLF_61_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_96 (.A(\b7_nYJ_BFM[261] ), .B(
        \b7_nYJ_BFM[134] ), .C(\b7_vFW_PlM[260] ), .D(
        \b7_vFW_PlM[133] ), .Y(b3_PLF_96_net_1));
    SLE \genblk9.b9_v_mzCDYXs[0]  (.D(b9_v_mzCDYXs_2), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[0] ));
    SLE \genblk9.b7_nYJ_BFM[79]  (.D(\b7_nYJ_BFM[78] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[79] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_10 (.A(\b7_nYJ_BFM[280] ), .B(
        \b7_nYJ_BFM[153] ), .C(\b7_vFW_PlM[279] ), .D(
        \b7_vFW_PlM[152] ), .Y(b3_PLF_10_net_1));
    SLE \genblk9.b7_nYJ_BFM[380]  (.D(\b7_nYJ_BFM[379] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[380] ));
    SLE \genblk9.b7_nYJ_BFM[308]  (.D(\b7_nYJ_BFM[307] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[308] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_s_9 (.A(VCC_net_1)
        , .B(\b12_2_St6KCa_jHv[9]_net_1 ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(un1_b12_2_St6KCa_jHv_cry_8_net_1), .S(
        un1_b12_2_St6KCa_jHv_s_9_S), .Y(), .FCO());
    SLE \genblk9.b7_nYJ_BFM[223]  (.D(\b7_nYJ_BFM[222] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[223] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_174 (.A(\b7_nYJ_BFM[377] ), .B(
        \b7_nYJ_BFM[121] ), .C(\b7_vFW_PlM[376] ), .D(
        \b7_vFW_PlM[120] ), .Y(b3_PLF_174_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[6]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNILNNS6_S[6] ), .Y(b9_v_mzCDYXs_6));
    SLE \genblk9.b7_nYJ_BFM[139]  (.D(\b7_nYJ_BFM[138] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[139] ));
    SLE \genblk9.b7_nYJ_BFM[114]  (.D(\b7_nYJ_BFM[113] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[114] ));
    SLE \genblk9.b7_nYJ_BFM[365]  (.D(\b7_nYJ_BFM[364] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[365] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_50 (.A(\b7_nYJ_BFM[195] ), .B(
        \b7_nYJ_BFM[68] ), .C(\b7_vFW_PlM[194] ), .D(\b7_vFW_PlM[67] ), 
        .Y(b3_PLF_50_net_1));
    SLE \genblk9.b7_nYJ_BFM[345]  (.D(\b7_nYJ_BFM[344] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[345] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_151 (.A(\b7_nYJ_BFM[345] ), .B(
        \b7_nYJ_BFM[89] ), .C(\b7_vFW_PlM[344] ), .D(\b7_vFW_PlM[88] ), 
        .Y(b3_PLF_151_net_1));
    SLE \genblk9.b7_nYJ_BFM[69]  (.D(\b7_nYJ_BFM[68] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[69] ));
    SLE \genblk9.b7_nYJ_BFM[122]  (.D(\b7_nYJ_BFM[121] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[122] ));
    SLE \b12_PSyi_KyDbLbb[9]  (.D(\b12_2_St6KCa_jHv[9]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[9]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[269]  (.D(\b7_nYJ_BFM[268] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[269] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_327 (.A(b3_PLF_180_net_1), .B(
        b3_PLF_179_net_1), .C(b3_PLF_178_net_1), .D(b3_PLF_177_net_1), 
        .Y(b3_PLF_327_net_1));
    SLE \genblk9.b7_nYJ_BFM[249]  (.D(\b7_nYJ_BFM[248] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[249] ));
    SLE \genblk9.b7_nYJ_BFM[185]  (.D(\b7_nYJ_BFM[184] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[185] ));
    SLE \genblk9.b7_nYJ_BFM[273]  (.D(\b7_nYJ_BFM[272] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[273] ));
    SLE \b8_FZFFLXYE[3]  (.D(\b12_2_St6KCa_jHv[3]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_181 (.A(\b7_nYJ_BFM[351] ), .B(
        \b7_nYJ_BFM[240] ), .C(\b7_vFW_PlM[350] ), .D(
        \b7_vFW_PlM[239] ), .Y(b3_PLF_181_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_120 (.A(\b7_nYJ_BFM[164] ), .B(
        \b7_nYJ_BFM[37] ), .C(\b7_vFW_PlM[163] ), .D(\b7_vFW_PlM[36] ), 
        .Y(b3_PLF_120_net_1));
    SLE \genblk9.b7_nYJ_BFM[183]  (.D(\b7_nYJ_BFM[182] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[183] ));
    SLE \genblk9.b7_nYJ_BFM[330]  (.D(\b7_nYJ_BFM[329] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[330] ));
    SLE \b8_FZFFLXYE[7]  (.D(\b12_2_St6KCa_jHv[7]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[7]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[172]  (.D(\b7_nYJ_BFM[171] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[172] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_13 (.A(\b7_nYJ_BFM[276] ), .B(
        \b7_nYJ_BFM[149] ), .C(\b7_vFW_PlM[275] ), .D(
        \b7_vFW_PlM[148] ), .Y(b3_PLF_13_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_123 (.A(\b7_nYJ_BFM[160] ), .B(
        \b7_nYJ_BFM[33] ), .C(\b7_vFW_PlM[159] ), .D(\b7_vFW_PlM[32] ), 
        .Y(b3_PLF_123_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_290 (.A(b3_PLF_32_net_1), .B(
        b3_PLF_31_net_1), .C(b3_PLF_30_net_1), .D(b3_PLF_29_net_1), .Y(
        b3_PLF_290_net_1));
    SLE \genblk9.b7_nYJ_BFM[292]  (.D(\b7_nYJ_BFM[291] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[292] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_87 (.A(\b7_nYJ_BFM[370] ), .B(
        \b7_nYJ_BFM[114] ), .C(\b7_vFW_PlM[369] ), .D(
        \b7_vFW_PlM[113] ), .Y(b3_PLF_87_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_39 (.A(\b7_nYJ_BFM[306] ), .B(
        \b7_nYJ_BFM[50] ), .C(\b7_vFW_PlM[305] ), .D(\b7_vFW_PlM[49] ), 
        .Y(b3_PLF_39_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_67 (.A(\b7_nYJ_BFM[268] ), .B(
        \b7_nYJ_BFM[157] ), .C(\b7_vFW_PlM[267] ), .D(
        \b7_vFW_PlM[156] ), .Y(b3_PLF_67_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_53 (.A(\b7_nYJ_BFM[175] ), .B(
        \b7_nYJ_BFM[64] ), .C(\b7_vFW_PlM[174] ), .D(\b7_vFW_PlM[63] ), 
        .Y(b3_PLF_53_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_144 (.A(\b7_nYJ_BFM[323] ), .B(
        \b7_nYJ_BFM[67] ), .C(\b7_vFW_PlM[322] ), .D(\b7_vFW_PlM[66] ), 
        .Y(b3_PLF_144_net_1));
    SLE \b12_2_St6KCa_jHv[4]  (.D(b12_2_St6KCa_jHv_3), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[4]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[78]  (.D(\b7_nYJ_BFM[77] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[78] ));
    SLE \genblk9.b7_nYJ_BFM[309]  (.D(\b7_nYJ_BFM[308] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[309] ));
    SLE \genblk9.b7_nYJ_BFM[135]  (.D(\b7_nYJ_BFM[134] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[135] ));
    SLE \genblk9.b7_nYJ_BFM[213]  (.D(\b7_nYJ_BFM[212] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[213] ));
    SLE \genblk9.b7_nYJ_BFM[184]  (.D(\b7_nYJ_BFM[183] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[184] ));
    SLE \genblk9.b7_nYJ_BFM[99]  (.D(\b7_nYJ_BFM[98] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[99] ));
    SLE \genblk9.b7_nYJ_BFM[133]  (.D(\b7_nYJ_BFM[132] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[133] ));
    SLE \genblk9.b7_nYJ_BFM[205]  (.D(\b7_nYJ_BFM[204] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[205] ));
    SLE \genblk9.b7_nYJ_BFM[112]  (.D(\b7_nYJ_BFM[111] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[112] ));
    SLE \genblk9.b7_nYJ_BFM[68]  (.D(\b7_nYJ_BFM[67] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[68] ));
    SLE \genblk9.b7_nYJ_BFM[43]  (.D(\b7_nYJ_BFM[42] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[43] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_26 (.A(\b7_nYJ_BFM[163] ), .B(
        \b7_nYJ_BFM[36] ), .C(\b7_vFW_PlM[162] ), .D(\b7_vFW_PlM[35] ), 
        .Y(b3_PLF_26_net_1));
    CFG4 #( .INIT(16'h8000) )  b8_jAA_KlCO_0_sqmuxa_6 (.A(
        \b12_2_St6KCa_jHv[9]_net_1 ), .B(\b12_2_St6KCa_jHv[2]_net_1 ), 
        .C(\b12_2_St6KCa_jHv[1]_net_1 ), .D(
        \b12_2_St6KCa_jHv[0]_net_1 ), .Y(b8_jAA_KlCO_0_sqmuxa_6_net_1));
    SLE \genblk9.b7_nYJ_BFM[86]  (.D(\b7_nYJ_BFM[85] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[86] ));
    SLE \b12_PSyi_KyDbLbb[6]  (.D(\b12_2_St6KCa_jHv[6]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_159 (.A(\b7_nYJ_BFM[174] ), .B(
        \b7_nYJ_BFM[63] ), .C(\b7_vFW_PlM[173] ), .D(\b7_vFW_PlM[62] ), 
        .Y(b3_PLF_159_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_84 (.A(\b7_nYJ_BFM[374] ), .B(
        \b7_nYJ_BFM[118] ), .C(\b7_vFW_PlM[373] ), .D(
        \b7_vFW_PlM[117] ), .Y(b3_PLF_84_net_1));
    SLE \genblk9.b7_nYJ_BFM[134]  (.D(\b7_nYJ_BFM[133] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[134] ));
    SLE \genblk9.b7_nYJ_BFM[157]  (.D(\b7_nYJ_BFM[156] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[157] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_7 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[7]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_6_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_7_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_7_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_64 (.A(\b7_nYJ_BFM[336] ), .B(
        \b7_nYJ_BFM[209] ), .C(\b7_vFW_PlM[335] ), .D(
        \b7_vFW_PlM[208] ), .Y(b3_PLF_64_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_359 (.A(b3_PLF_308_net_1), .B(
        b3_PLF_307_net_1), .C(b3_PLF_306_net_1), .D(b3_PLF_305_net_1), 
        .Y(b3_PLF_359_net_1));
    SLE \genblk9.b7_nYJ_BFM[101]  (.D(\b7_nYJ_BFM[100] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[101] ));
    SLE \genblk9.b7_nYJ_BFM[1]  (.D(\b7_nYJ_BFM[0] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[1] ));
    SLE \genblk9.b7_nYJ_BFM[366]  (.D(\b7_nYJ_BFM[365] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[366] ));
    SLE \genblk9.b7_nYJ_BFM[128]  (.D(\b7_nYJ_BFM[127] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[128] ));
    SLE \genblk9.b7_nYJ_BFM[346]  (.D(\b7_nYJ_BFM[345] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[346] ));
    SLE \genblk9.b7_nYJ_BFM[283]  (.D(\b7_nYJ_BFM[282] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[283] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_95 (.A(\b7_nYJ_BFM[263] ), .B(
        \b7_nYJ_BFM[7] ), .C(\b7_vFW_PlM[262] ), .D(\b7_vFW_PlM[6] ), 
        .Y(b3_PLF_95_net_1));
    SLE \genblk9.b7_nYJ_BFM[55]  (.D(\b7_nYJ_BFM[54] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[55] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_356 (.A(b3_PLF_296_net_1), .B(
        b3_PLF_295_net_1), .C(b3_PLF_294_net_1), .D(b3_PLF_293_net_1), 
        .Y(b3_PLF_356_net_1));
    SLE \genblk9.b7_nYJ_BFM[291]  (.D(\b7_nYJ_BFM[290] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[291] ));
    SLE \genblk9.b7_nYJ_BFM[357]  (.D(\b7_nYJ_BFM[356] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[357] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_318 (.A(b3_PLF_144_net_1), .B(
        b3_PLF_143_net_1), .C(b3_PLF_142_net_1), .D(b3_PLF_141_net_1), 
        .Y(b3_PLF_318_net_1));
    SLE \genblk9.b7_nYJ_BFM[98]  (.D(\b7_nYJ_BFM[97] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[98] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_98 (.A(\b7_nYJ_BFM[259] ), .B(
        \b7_nYJ_BFM[3] ), .C(\b7_vFW_PlM[258] ), .D(\b7_vFW_PlM[2] ), 
        .Y(b3_PLF_98_net_1));
    SLE \genblk9.b7_nYJ_BFM[182]  (.D(\b7_nYJ_BFM[181] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[182] ));
    SLE \genblk9.b7_nYJ_BFM[260]  (.D(\b7_nYJ_BFM[259] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[260] ));
    CFG2 #( .INIT(4'h8) )  N_850_a2_1 (.A(b10_OFWNT9khFt), .B(
        IICE_comm2iice_10), .Y(N_850_a2_1_net_1));
    SLE \genblk9.b7_nYJ_BFM[35]  (.D(\b7_nYJ_BFM[34] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[35] ));
    SLE \genblk9.b7_nYJ_BFM[240]  (.D(\b7_nYJ_BFM[239] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[240] ));
    SLE \genblk9.b7_nYJ_BFM[44]  (.D(\b7_nYJ_BFM[43] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[44] ));
    SLE \genblk9.b7_nYJ_BFM[358]  (.D(\b7_nYJ_BFM[357] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[358] ));
    SLE \genblk9.b7_nYJ_BFM[178]  (.D(\b7_nYJ_BFM[177] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[178] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_298 (.A(b3_PLF_64_net_1), .B(
        b3_PLF_63_net_1), .C(b3_PLF_62_net_1), .D(b3_PLF_61_net_1), .Y(
        b3_PLF_298_net_1));
    SLE \genblk9.b7_nYJ_BFM[22]  (.D(\b7_nYJ_BFM[21] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[22] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_41 (.A(\b7_nYJ_BFM[159] ), .B(
        \b7_nYJ_BFM[48] ), .C(\b7_vFW_PlM[158] ), .D(\b7_vFW_PlM[47] ), 
        .Y(b3_PLF_41_net_1));
    CFG2 #( .INIT(4'hE) )  b8_jAA_KlCO_RNO (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .Y(
        b8_jAA_KlCO_RNO_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_314 (.A(b3_PLF_128_net_1), .B(
        b3_PLF_127_net_1), .C(b3_PLF_126_net_1), .D(b3_PLF_125_net_1), 
        .Y(b3_PLF_314_net_1));
    SLE \genblk9.b7_nYJ_BFM[233]  (.D(\b7_nYJ_BFM[232] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[233] ));
    SLE \genblk9.b7_nYJ_BFM[364]  (.D(\b7_nYJ_BFM[363] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[364] ));
    SLE \genblk9.b7_nYJ_BFM[344]  (.D(\b7_nYJ_BFM[343] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[344] ));
    SLE \b8_FZFFLXYE[6]  (.D(\b12_2_St6KCa_jHv[6]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[6]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[132]  (.D(\b7_nYJ_BFM[131] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[132] ));
    SLE \b12_PSyi_KyDbLbb[1]  (.D(\b12_2_St6KCa_jHv[1]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_0 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[0]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_s_0_532_FCO), .S(
        un1_b12_2_St6KCa_jHv_cry_0_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_0_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_301 (.A(b3_PLF_76_net_1), .B(
        b3_PLF_75_net_1), .C(b3_PLF_74_net_1), .D(b3_PLF_73_net_1), .Y(
        b3_PLF_301_net_1));
    SLE \genblk9.b7_nYJ_BFM[106]  (.D(\b7_nYJ_BFM[105] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[106] ));
    SLE \genblk9.b7_nYJ_BFM[118]  (.D(\b7_nYJ_BFM[117] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[118] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_312 (.A(b3_PLF_120_net_1), .B(
        b3_PLF_119_net_1), .C(b3_PLF_118_net_1), .D(b3_PLF_117_net_1), 
        .Y(b3_PLF_312_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_305 (.A(b3_PLF_92_net_1), .B(
        b3_PLF_91_net_1), .C(b3_PLF_90_net_1), .D(b3_PLF_89_net_1), .Y(
        b3_PLF_305_net_1));
    SLE \genblk9.b7_nYJ_BFM[4]  (.D(\b7_nYJ_BFM[3] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[4] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_12 (.A(\b7_nYJ_BFM[278] ), .B(
        \b7_nYJ_BFM[22] ), .C(\b7_vFW_PlM[277] ), .D(\b7_vFW_PlM[21] ), 
        .Y(b3_PLF_12_net_1));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b9_v_mzCDYXs_RNIRFPF3[7]  (.A(
        \b9_v_mzCDYXs[9] ), .B(\b9_v_mzCDYXs[7] ), .C(m9_e_6), .D(
        m9_e_5), .Y(N_24_mux));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_167 (.A(\b7_nYJ_BFM[355] ), .B(
        \b7_nYJ_BFM[99] ), .C(\b7_vFW_PlM[354] ), .D(\b7_vFW_PlM[98] ), 
        .Y(b3_PLF_167_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_106 (.A(\b7_nYJ_BFM[279] ), .B(
        \b7_nYJ_BFM[152] ), .C(\b7_vFW_PlM[278] ), .D(
        \b7_vFW_PlM[151] ), .Y(b3_PLF_106_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_1 (.A(\b7_nYJ_BFM[260] ), .B(
        \b7_nYJ_BFM[133] ), .C(\b7_vFW_PlM[259] ), .D(
        \b7_vFW_PlM[132] ), .Y(b3_PLF_1_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_52 (.A(\b7_nYJ_BFM[320] ), .B(
        \b7_nYJ_BFM[193] ), .C(\b7_vFW_PlM[319] ), .D(
        \b7_vFW_PlM[192] ), .Y(b3_PLF_52_net_1));
    SLE \genblk9.b7_nYJ_BFM[359]  (.D(\b7_nYJ_BFM[358] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[359] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[9]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_s_9_S), .Y(b12_2_St6KCa_jHv_8));
    SLE \genblk9.b7_nYJ_BFM[51]  (.D(\b7_nYJ_BFM[50] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[51] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_25 (.A(\b7_nYJ_BFM[292] ), .B(
        \b7_nYJ_BFM[165] ), .C(\b7_vFW_PlM[291] ), .D(
        \b7_vFW_PlM[164] ), .Y(b3_PLF_25_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_47 (.A(\b7_nYJ_BFM[199] ), .B(
        \b7_nYJ_BFM[72] ), .C(\b7_vFW_PlM[198] ), .D(\b7_vFW_PlM[71] ), 
        .Y(b3_PLF_47_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_118 (.A(\b7_nYJ_BFM[295] ), .B(
        \b7_nYJ_BFM[39] ), .C(\b7_vFW_PlM[294] ), .D(\b7_vFW_PlM[38] ), 
        .Y(b3_PLF_118_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_5 (.A(\b7_nYJ_BFM[367] ), .B(
        \b7_nYJ_BFM[111] ), .C(\b7_vFW_PlM[366] ), .D(
        \b7_vFW_PlM[110] ), .Y(b3_PLF_5_net_1));
    SLE \genblk9.b7_nYJ_BFM[255]  (.D(\b7_nYJ_BFM[254] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[255] ));
    SLE \b12_PSyi_KyDbLbb[4]  (.D(\b12_2_St6KCa_jHv[4]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[4]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[31]  (.D(\b7_nYJ_BFM[30] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[31] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_36 (.A(\b7_nYJ_BFM[310] ), .B(
        \b7_nYJ_BFM[54] ), .C(\b7_vFW_PlM[309] ), .D(\b7_vFW_PlM[53] ), 
        .Y(b3_PLF_36_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_28 (.A(\b7_nYJ_BFM[288] ), .B(
        \b7_nYJ_BFM[161] ), .C(\b7_vFW_PlM[287] ), .D(
        \b7_vFW_PlM[160] ), .Y(b3_PLF_28_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_162 (.A(\b7_nYJ_BFM[361] ), .B(
        \b7_nYJ_BFM[234] ), .C(\b7_vFW_PlM[360] ), .D(
        \b7_vFW_PlM[233] ), .Y(b3_PLF_162_net_1));
    SLE \genblk9.b7_nYJ_BFM[3]  (.D(\b7_nYJ_BFM[2] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[3] ));
    SLE \genblk9.b7_nYJ_BFM[10]  (.D(\b7_nYJ_BFM[9] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[10] ));
    SLE \genblk9.b7_nYJ_BFM[222]  (.D(\b7_nYJ_BFM[221] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[222] ));
    SLE \genblk9.b7_nYJ_BFM[296]  (.D(\b7_nYJ_BFM[295] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[296] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_136 (.A(\b7_nYJ_BFM[142] ), .B(
        \b7_nYJ_BFM[31] ), .C(\b7_vFW_PlM[141] ), .D(\b7_vFW_PlM[30] ), 
        .Y(b3_PLF_136_net_1));
    SLE \genblk9.b7_nYJ_BFM[188]  (.D(\b7_nYJ_BFM[187] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[188] ));
    CFG3 #( .INIT(8'hE2) )  b7_yYh03wy_u_0_m2 (.A(b4_ycsM), .B(
        IICE_comm2iice_5), .C(ttdo), .Y(b7_yYh03wy_u_0_m2_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_71 (.A(\b7_nYJ_BFM[231] ), .B(
        \b7_nYJ_BFM[104] ), .C(\b7_vFW_PlM[230] ), .D(
        \b7_vFW_PlM[103] ), .Y(b3_PLF_71_net_1));
    SLE \b12_2_St6KCa_jHv[3]  (.D(b12_2_St6KCa_jHv_2), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_105 (.A(\b7_nYJ_BFM[281] ), .B(
        \b7_nYJ_BFM[25] ), .C(\b7_vFW_PlM[280] ), .D(\b7_vFW_PlM[24] ), 
        .Y(b3_PLF_105_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_372 (.A(b3_PLF_360_net_1), .B(
        b3_PLF_359_net_1), .C(b3_PLF_358_net_1), .D(b3_PLF_357_net_1), 
        .Y(b3_PLF_372_net_1));
    SLE \b12_PSyi_KyDbLbb[2]  (.D(\b12_2_St6KCa_jHv[2]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[2]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[151]  (.D(\b7_nYJ_BFM[150] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[151] ));
    SLE \genblk9.b7_nYJ_BFM[362]  (.D(\b7_nYJ_BFM[361] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[362] ));
    SLE \genblk9.b7_nYJ_BFM[342]  (.D(\b7_nYJ_BFM[341] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[342] ));
    SLE \genblk9.b7_nYJ_BFM[272]  (.D(\b7_nYJ_BFM[271] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[272] ));
    SLE \genblk9.b7_nYJ_BFM[87]  (.D(\b7_nYJ_BFM[86] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[87] ));
    SLE \genblk9.b7_nYJ_BFM[361]  (.D(\b7_nYJ_BFM[360] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[361] ));
    ARI1 #( .INIT(20'h40040) )  \genblk9.b7_nYJ_BFM_RNIJQFE4[383]  (.A(
        b8_SoWGfWYY), .B(N_24_mux), .C(N_850_a2_1_net_1), .D(
        b8_nYJ_TqLY), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        b9_v_mzCDYXs_cry_0_cy));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[0]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNIUDLP4_S[0] ), .Y(b9_v_mzCDYXs_2));
    SLE \genblk9.b7_nYJ_BFM[341]  (.D(\b7_nYJ_BFM[340] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[341] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_44 (.A(\b7_nYJ_BFM[347] ), .B(
        \b7_nYJ_BFM[219] ), .C(\b7_vFW_PlM[346] ), .D(
        \b7_vFW_PlM[218] ), .Y(b3_PLF_44_net_1));
    SLE \genblk9.b7_nYJ_BFM[267]  (.D(\b7_nYJ_BFM[266] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[267] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_291 (.A(b3_PLF_36_net_1), .B(
        b3_PLF_35_net_1), .C(b3_PLF_34_net_1), .D(b3_PLF_33_net_1), .Y(
        b3_PLF_291_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIA2R45[1]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[1] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_0), .S(\b9_v_mzCDYXs_RNIA2R45_S[1] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_1));
    SLE \genblk9.b7_nYJ_BFM[247]  (.D(\b7_nYJ_BFM[246] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[247] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_296 (.A(b3_PLF_56_net_1), .B(
        b3_PLF_55_net_1), .C(b3_PLF_54_net_1), .D(b3_PLF_53_net_1), .Y(
        b3_PLF_296_net_1));
    SLE \genblk9.b7_nYJ_BFM[138]  (.D(\b7_nYJ_BFM[137] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[138] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_178 (.A(\b7_nYJ_BFM[371] ), .B(
        \b7_nYJ_BFM[244] ), .C(\b7_vFW_PlM[370] ), .D(
        \b7_vFW_PlM[243] ), .Y(b3_PLF_178_net_1));
    SLE \genblk9.b7_nYJ_BFM[6]  (.D(\b7_nYJ_BFM[5] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[6] ));
    SLE \genblk9.b7_nYJ_BFM[29]  (.D(\b7_nYJ_BFM[28] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[29] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_135 (.A(\b7_nYJ_BFM[287] ), .B(
        \b7_nYJ_BFM[176] ), .C(\b7_vFW_PlM[286] ), .D(
        \b7_vFW_PlM[175] ), .Y(b3_PLF_135_net_1));
    SLE \genblk9.b7_nYJ_BFM[212]  (.D(\b7_nYJ_BFM[211] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[212] ));
    SLE \genblk9.b9_v_mzCDYXs[5]  (.D(b9_v_mzCDYXs_7), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[5] ));
    b19_nczQ_DYg_YFaRM_oUoP_24s_1s_x_0 samplerStatus (
        .b12_PSyi_KyDbLbb({\b12_PSyi_KyDbLbb[9]_net_1 , 
        \b12_PSyi_KyDbLbb[8]_net_1 , \b12_PSyi_KyDbLbb[7]_net_1 , 
        \b12_PSyi_KyDbLbb[6]_net_1 , \b12_PSyi_KyDbLbb[5]_net_1 , 
        \b12_PSyi_KyDbLbb[4]_net_1 , \b12_PSyi_KyDbLbb[3]_net_1 , 
        \b12_PSyi_KyDbLbb[2]_net_1 , \b12_PSyi_KyDbLbb[1]_net_1 , 
        \b12_PSyi_KyDbLbb[0]_net_1 }), .b8_FZFFLXYE({
        \b8_FZFFLXYE[9]_net_1 , \b8_FZFFLXYE[8]_net_1 , 
        \b8_FZFFLXYE[7]_net_1 , \b8_FZFFLXYE[6]_net_1 , 
        \b8_FZFFLXYE[5]_net_1 , \b8_FZFFLXYE[4]_net_1 , 
        \b8_FZFFLXYE[3]_net_1 , \b8_FZFFLXYE[2]_net_1 , 
        \b8_FZFFLXYE[1]_net_1 , \b8_FZFFLXYE[0]_net_1 }), 
        .IICE_comm2iice_6(IICE_comm2iice_11), .IICE_comm2iice_4(
        IICE_comm2iice_9), .IICE_comm2iice_5(IICE_comm2iice_10), 
        .IICE_comm2iice_0(IICE_comm2iice_5), .IICE_comm2iice_1(
        IICE_comm2iice_6), .ttdo(ttdo), .un1_b5_OvyH3(un1_b5_OvyH3), 
        .b8_jAA_KlCO(b8_jAA_KlCO_net_1), .N_21(N_21));
    SLE \genblk9.b7_nYJ_BFM[46]  (.D(\b7_nYJ_BFM[45] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[46] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_77 (.A(\b7_nYJ_BFM[207] ), .B(
        \b7_nYJ_BFM[96] ), .C(\b7_vFW_PlM[206] ), .D(\b7_vFW_PlM[95] ), 
        .Y(b3_PLF_77_net_1));
    SLE \genblk9.b7_nYJ_BFM[221]  (.D(\b7_nYJ_BFM[220] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[221] ));
    SLE \genblk9.b7_nYJ_BFM[160]  (.D(\b7_nYJ_BFM[159] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[160] ));
    SLE \genblk9.b7_nYJ_BFM[140]  (.D(\b7_nYJ_BFM[139] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[140] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_310 (.A(b3_PLF_112_net_1), .B(
        b3_PLF_111_net_1), .C(b3_PLF_110_net_1), .D(b3_PLF_109_net_1), 
        .Y(b3_PLF_310_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_157 (.A(\b7_nYJ_BFM[337] ), .B(
        \b7_nYJ_BFM[81] ), .C(\b7_vFW_PlM[336] ), .D(\b7_vFW_PlM[80] ), 
        .Y(b3_PLF_157_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_101 (.A(\b7_nYJ_BFM[350] ), .B(
        \b7_nYJ_BFM[239] ), .C(\b7_vFW_PlM[349] ), .D(
        \b7_vFW_PlM[238] ), .Y(b3_PLF_101_net_1));
    SLE \b12_2_St6KCa_jHv[9]  (.D(b12_2_St6KCa_jHv_8), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[9]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[156]  (.D(\b7_nYJ_BFM[155] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[156] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_4 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[4]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_3_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_4_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_4_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_148 (.A(\b7_nYJ_BFM[269] ), .B(
        \b7_nYJ_BFM[158] ), .C(\b7_vFW_PlM[268] ), .D(
        \b7_vFW_PlM[157] ), .Y(b3_PLF_148_net_1));
    SLE \genblk9.b7_nYJ_BFM[271]  (.D(\b7_nYJ_BFM[270] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[271] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_187 (.A(\b7_nYJ_BFM[264] ), .B(
        \b7_nYJ_BFM[8] ), .C(\b7_vFW_PlM[263] ), .D(\b7_vFW_PlM[7] ), 
        .Y(b3_PLF_187_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_89 (.A(\b7_nYJ_BFM[223] ), .B(
        \b7_nYJ_BFM[112] ), .C(\b7_vFW_PlM[222] ), .D(
        \b7_vFW_PlM[111] ), .Y(b3_PLF_89_net_1));
    SLE \genblk9.b7_nYJ_BFM[305]  (.D(\b7_nYJ_BFM[304] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[305] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_69 (.A(\b7_nYJ_BFM[106] ), .B(
        \b7_nYJ_BFM[11] ), .C(\b7_vFW_PlM[105] ), .D(\b7_vFW_PlM[10] ), 
        .Y(b3_PLF_69_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_313 (.A(b3_PLF_124_net_1), .B(
        b3_PLF_123_net_1), .C(b3_PLF_122_net_1), .D(b3_PLF_121_net_1), 
        .Y(b3_PLF_313_net_1));
    SLE \genblk9.b7_nYJ_BFM[28]  (.D(\b7_nYJ_BFM[27] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[28] ));
    CFG2 #( .INIT(4'h8) )  b8_jAA_KlCO_0_sqmuxa_4 (.A(
        \b12_2_St6KCa_jHv[5]_net_1 ), .B(\b12_2_St6KCa_jHv[6]_net_1 ), 
        .Y(b8_jAA_KlCO_0_sqmuxa_4_net_1));
    SLE \genblk9.b7_nYJ_BFM[282]  (.D(\b7_nYJ_BFM[281] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[282] ));
    SLE \genblk9.b7_nYJ_BFM[70]  (.D(\b7_nYJ_BFM[69] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[70] ));
    SLE \genblk9.b7_nYJ_BFM[209]  (.D(\b7_nYJ_BFM[208] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[209] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_35 (.A(\b7_nYJ_BFM[183] ), .B(
        \b7_nYJ_BFM[56] ), .C(\b7_vFW_PlM[182] ), .D(\b7_vFW_PlM[55] ), 
        .Y(b3_PLF_35_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_152 (.A(\b7_nYJ_BFM[343] ), .B(
        \b7_nYJ_BFM[216] ), .C(\b7_vFW_PlM[342] ), .D(
        \b7_vFW_PlM[215] ), .Y(b3_PLF_152_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_74 (.A(\b7_nYJ_BFM[227] ), .B(
        \b7_nYJ_BFM[100] ), .C(\b7_vFW_PlM[226] ), .D(\b7_vFW_PlM[99] )
        , .Y(b3_PLF_74_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_321 (.A(b3_PLF_156_net_1), .B(
        b3_PLF_155_net_1), .C(b3_PLF_154_net_1), .D(b3_PLF_153_net_1), 
        .Y(b3_PLF_321_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_38 (.A(\b7_nYJ_BFM[179] ), .B(
        \b7_nYJ_BFM[52] ), .C(\b7_vFW_PlM[178] ), .D(\b7_vFW_PlM[51] ), 
        .Y(b3_PLF_38_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_131 (.A(\b7_nYJ_BFM[309] ), .B(
        \b7_nYJ_BFM[53] ), .C(\b7_vFW_PlM[308] ), .D(\b7_vFW_PlM[52] ), 
        .Y(b3_PLF_131_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_182 (.A(\b7_nYJ_BFM[206] ), .B(
        \b7_nYJ_BFM[95] ), .C(\b7_vFW_PlM[205] ), .D(\b7_vFW_PlM[94] ), 
        .Y(b3_PLF_182_net_1));
    SLE \genblk9.b7_nYJ_BFM[211]  (.D(\b7_nYJ_BFM[210] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[211] ));
    SLE \genblk9.b7_nYJ_BFM[60]  (.D(\b7_nYJ_BFM[59] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[60] ));
    SLE \genblk9.b7_nYJ_BFM[323]  (.D(\b7_nYJ_BFM[322] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[323] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_325 (.A(b3_PLF_172_net_1), .B(
        b3_PLF_171_net_1), .C(b3_PLF_170_net_1), .D(b3_PLF_169_net_1), 
        .Y(b3_PLF_325_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_126 (.A(\b7_nYJ_BFM[348] ), .B(
        \b7_nYJ_BFM[92] ), .C(\b7_vFW_PlM[347] ), .D(\b7_vFW_PlM[91] ), 
        .Y(b3_PLF_126_net_1));
    SLE \genblk9.b7_nYJ_BFM[232]  (.D(\b7_nYJ_BFM[231] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[232] ));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b9_v_mzCDYXs_RNI24NC1[3]  (.A(
        \b9_v_mzCDYXs[8] ), .B(\b9_v_mzCDYXs[6] ), .C(
        \b9_v_mzCDYXs[5] ), .D(\b9_v_mzCDYXs[3] ), .Y(m9_e_6));
    SLE \genblk9.b7_nYJ_BFM[373]  (.D(\b7_nYJ_BFM[372] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[373] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_109 (.A(\b7_nYJ_BFM[275] ), .B(
        \b7_nYJ_BFM[148] ), .C(\b7_vFW_PlM[274] ), .D(
        \b7_vFW_PlM[147] ), .Y(b3_PLF_109_net_1));
    SLE \b12_2_St6KCa_jHv[8]  (.D(b12_2_St6KCa_jHv_7), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[8]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[13]  (.D(\b7_nYJ_BFM[12] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[13] ));
    SLE \genblk9.b9_v_mzCDYXs[9]  (.D(b9_v_mzCDYXs_3), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[9] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_373 (.A(b3_PLF_364_net_1), .B(
        b3_PLF_363_net_1), .C(b3_PLF_362_net_1), .D(b3_PLF_361_net_1), 
        .Y(b3_PLF_373_net_1));
    SLE \genblk9.b7_nYJ_BFM[226]  (.D(\b7_nYJ_BFM[225] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[226] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_309 (.A(b3_PLF_108_net_1), .B(
        b3_PLF_107_net_1), .C(b3_PLF_106_net_1), .D(b3_PLF_105_net_1), 
        .Y(b3_PLF_309_net_1));
    SLE \b12_PSyi_KyDbLbb[0]  (.D(\b12_2_St6KCa_jHv[0]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[0]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[197]  (.D(\b7_nYJ_BFM[196] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[197] ));
    SLE \genblk9.b7_nYJ_BFM[90]  (.D(\b7_nYJ_BFM[89] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[90] ));
    SLE \genblk9.b7_nYJ_BFM[264]  (.D(\b7_nYJ_BFM[263] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[264] ));
    SLE \genblk9.b7_nYJ_BFM[52]  (.D(\b7_nYJ_BFM[51] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[52] ));
    SLE \genblk9.b7_nYJ_BFM[244]  (.D(\b7_nYJ_BFM[243] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[244] ));
    SLE \genblk9.b7_nYJ_BFM[281]  (.D(\b7_nYJ_BFM[280] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[281] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_90 (.A(\b7_nYJ_BFM[334] ), .B(
        \b7_nYJ_BFM[78] ), .C(\b7_vFW_PlM[333] ), .D(\b7_vFW_PlM[77] ), 
        .Y(b3_PLF_90_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_306 (.A(b3_PLF_96_net_1), .B(
        b3_PLF_95_net_1), .C(b3_PLF_94_net_1), .D(b3_PLF_93_net_1), .Y(
        b3_PLF_306_net_1));
    SLE \genblk9.b7_nYJ_BFM[313]  (.D(\b7_nYJ_BFM[312] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[313] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_125 (.A(\b7_nYJ_BFM[237] ), .B(
        \b7_nYJ_BFM[126] ), .C(\b7_vFW_PlM[236] ), .D(
        \b7_vFW_PlM[125] ), .Y(b3_PLF_125_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[5]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNI4UHH6_S[5] ), .Y(b9_v_mzCDYXs_7));
    SLE \genblk9.b7_nYJ_BFM[276]  (.D(\b7_nYJ_BFM[275] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[276] ));
    SLE \genblk9.b7_nYJ_BFM[32]  (.D(\b7_nYJ_BFM[31] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[32] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_139 (.A(\b7_nYJ_BFM[329] ), .B(
        \b7_nYJ_BFM[202] ), .C(\b7_vFW_PlM[328] ), .D(
        \b7_vFW_PlM[201] ), .Y(b3_PLF_139_net_1));
    SLE \genblk9.b7_nYJ_BFM[268]  (.D(\b7_nYJ_BFM[267] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[268] ));
    SLE \genblk9.b7_nYJ_BFM[248]  (.D(\b7_nYJ_BFM[247] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[248] ));
    SLE \genblk9.b7_nYJ_BFM[306]  (.D(\b7_nYJ_BFM[305] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[306] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_288 (.A(b3_PLF_24_net_1), .B(
        b3_PLF_23_net_1), .C(b3_PLF_22_net_1), .D(b3_PLF_21_net_1), .Y(
        b3_PLF_288_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_317 (.A(b3_PLF_140_net_1), .B(
        b3_PLF_139_net_1), .C(b3_PLF_138_net_1), .D(b3_PLF_137_net_1), 
        .Y(b3_PLF_317_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_164 (.A(\b7_nYJ_BFM[359] ), .B(
        \b7_nYJ_BFM[103] ), .C(\b7_vFW_PlM[358] ), .D(
        \b7_vFW_PlM[102] ), .Y(b3_PLF_164_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_294 (.A(b3_PLF_48_net_1), .B(
        b3_PLF_47_net_1), .C(b3_PLF_46_net_1), .D(b3_PLF_45_net_1), .Y(
        b3_PLF_294_net_1));
    SLE \genblk9.b7_nYJ_BFM[231]  (.D(\b7_nYJ_BFM[230] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[231] ));
    SLE \genblk9.b7_nYJ_BFM[14]  (.D(\b7_nYJ_BFM[13] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[14] ));
    SLE \genblk9.b7_nYJ_BFM[169]  (.D(\b7_nYJ_BFM[168] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[169] ));
    SLE \genblk9.b7_nYJ_BFM[200]  (.D(\b7_nYJ_BFM[199] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[200] ));
    SLE \genblk9.b7_nYJ_BFM[149]  (.D(\b7_nYJ_BFM[148] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[149] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_110 (.A(\b7_nYJ_BFM[146] ), .B(
        \b7_nYJ_BFM[19] ), .C(\b7_vFW_PlM[145] ), .D(\b7_vFW_PlM[18] ), 
        .Y(b3_PLF_110_net_1));
    SLE \genblk9.b7_nYJ_BFM[7]  (.D(\b7_nYJ_BFM[6] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[7] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_93 (.A(\b7_nYJ_BFM[265] ), .B(
        \b7_nYJ_BFM[138] ), .C(\b7_vFW_PlM[264] ), .D(
        \b7_vFW_PlM[137] ), .Y(b3_PLF_93_net_1));
    SLE \genblk9.b7_nYJ_BFM[47]  (.D(\b7_nYJ_BFM[46] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[47] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_6 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[6]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_5_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_6_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_6_net_1));
    SLE \genblk9.b7_nYJ_BFM[216]  (.D(\b7_nYJ_BFM[215] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[216] ));
    SLE \genblk9.b7_nYJ_BFM[85]  (.D(\b7_nYJ_BFM[84] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[85] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_113 (.A(\b7_nYJ_BFM[110] ), .B(
        \b7_nYJ_BFM[15] ), .C(\b7_vFW_PlM[109] ), .D(\b7_vFW_PlM[14] ), 
        .Y(b3_PLF_113_net_1));
    SLE \genblk9.b7_nYJ_BFM[0]  (.D(b8_nYJ_TqLY), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(VCC_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[0] ));
    SLE \genblk9.b7_nYJ_BFM[355]  (.D(\b7_nYJ_BFM[354] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[355] ));
    SLE \genblk9.b7_nYJ_BFM[383]  (.D(\b7_nYJ_BFM[382] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b8_nYJ_TqLY));
    SLE \genblk9.b7_nYJ_BFM[360]  (.D(\b7_nYJ_BFM[359] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[360] ));
    SLE \genblk9.b7_nYJ_BFM[304]  (.D(\b7_nYJ_BFM[303] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[304] ));
    SLE \genblk9.b7_nYJ_BFM[259]  (.D(\b7_nYJ_BFM[258] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[259] ));
    SLE \genblk9.b7_nYJ_BFM[340]  (.D(\b7_nYJ_BFM[339] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[340] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_49 (.A(\b7_nYJ_BFM[324] ), .B(
        \b7_nYJ_BFM[197] ), .C(\b7_vFW_PlM[323] ), .D(
        \b7_vFW_PlM[196] ), .Y(b3_PLF_49_net_1));
    CFG4 #( .INIT(16'h0020) )  b12_PSyi_KyDbLbb_0_sqmuxa (.A(
        b11_PSyil9s_FMZ), .B(b9_PSyil9s_2_net_1), .C(b4_2o_z), .D(
        b8_SoWGfWYY), .Y(b12_PSyi_KyDbLbb_0_sqmuxa_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_86 (.A(\b7_nYJ_BFM[243] ), .B(
        \b7_nYJ_BFM[116] ), .C(\b7_vFW_PlM[242] ), .D(
        \b7_vFW_PlM[115] ), .Y(b3_PLF_86_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_121 (.A(\b7_nYJ_BFM[291] ), .B(
        \b7_nYJ_BFM[35] ), .C(\b7_vFW_PlM[290] ), .D(\b7_vFW_PlM[34] ), 
        .Y(b3_PLF_121_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[1]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_1_S), .Y(b12_2_St6KCa_jHv_0));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[7]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_7_S), .Y(b12_2_St6KCa_jHv_6));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_66 (.A(\b7_nYJ_BFM[302] ), .B(
        \b7_nYJ_BFM[46] ), .C(\b7_vFW_PlM[301] ), .D(\b7_vFW_PlM[45] ), 
        .Y(b3_PLF_66_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_20 (.A(\b7_nYJ_BFM[315] ), .B(
        \b7_nYJ_BFM[187] ), .C(\b7_vFW_PlM[314] ), .D(
        \b7_vFW_PlM[186] ), .Y(b3_PLF_20_net_1));
    SLE \genblk9.b7_nYJ_BFM[165]  (.D(\b7_nYJ_BFM[164] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[165] ));
    SLE \genblk9.b7_nYJ_BFM[145]  (.D(\b7_nYJ_BFM[144] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[145] ));
    SLE \genblk9.b7_nYJ_BFM[73]  (.D(\b7_nYJ_BFM[72] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[73] ));
    SLE \genblk9.b7_nYJ_BFM[333]  (.D(\b7_nYJ_BFM[332] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[333] ));
    SLE \genblk9.b7_nYJ_BFM[163]  (.D(\b7_nYJ_BFM[162] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[163] ));
    SLE \genblk9.b7_nYJ_BFM[295]  (.D(\b7_nYJ_BFM[294] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[295] ));
    SLE \genblk9.b7_nYJ_BFM[143]  (.D(\b7_nYJ_BFM[142] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[143] ));
    SLE \genblk9.b7_nYJ_BFM[286]  (.D(\b7_nYJ_BFM[285] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[286] ));
    SLE \genblk9.b7_nYJ_BFM[5]  (.D(\b7_nYJ_BFM[4] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[5] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_170 (.A(\b7_nYJ_BFM[335] ), .B(
        \b7_nYJ_BFM[79] ), .C(\b7_vFW_PlM[334] ), .D(\b7_vFW_PlM[78] ), 
        .Y(b3_PLF_170_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_173 (.A(\b7_nYJ_BFM[250] ), .B(
        \b7_nYJ_BFM[139] ), .C(\b7_vFW_PlM[249] ), .D(
        \b7_vFW_PlM[138] ), .Y(b3_PLF_173_net_1));
    SLE \genblk9.b7_nYJ_BFM[63]  (.D(\b7_nYJ_BFM[62] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[63] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_0 (.A(\b7_nYJ_BFM[262] ), .B(
        \b7_nYJ_BFM[6] ), .C(\b7_vFW_PlM[261] ), .D(\b7_vFW_PlM[5] ), 
        .Y(b3_PLF_0_net_1));
    SLE \genblk9.b7_nYJ_BFM[81]  (.D(\b7_nYJ_BFM[80] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[81] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_23 (.A(\b7_nYJ_BFM[167] ), .B(
        \b7_nYJ_BFM[40] ), .C(\b7_vFW_PlM[166] ), .D(\b7_vFW_PlM[39] ), 
        .Y(b3_PLF_23_net_1));
    SLE \genblk9.b7_nYJ_BFM[164]  (.D(\b7_nYJ_BFM[163] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[164] ));
    SLE \genblk9.b7_nYJ_BFM[2]  (.D(\b7_nYJ_BFM[1] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[2] ));
    SLE \genblk9.b7_nYJ_BFM[144]  (.D(\b7_nYJ_BFM[143] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[144] ));
    SLE \genblk9.b7_nYJ_BFM[59]  (.D(\b7_nYJ_BFM[58] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[59] ));
    SLE \genblk9.b7_nYJ_BFM[191]  (.D(\b7_nYJ_BFM[190] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[191] ));
    SLE \genblk9.b7_nYJ_BFM[236]  (.D(\b7_nYJ_BFM[235] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[236] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_3 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[3]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_2_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_3_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_3_net_1));
    CFG4 #( .INIT(16'hFEEE) )  b3_PLF_281 (.A(\un1_b4_BVmQ[265] ), .B(
        b3_PLF_186_net_1), .C(\b7_nYJ_BFM[155] ), .D(\b7_vFW_PlM[154] )
        , .Y(b3_PLF_281_net_1));
    SLE \genblk9.b7_nYJ_BFM[39]  (.D(\b7_nYJ_BFM[38] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[39] ));
    SLE \genblk9.b7_nYJ_BFM[302]  (.D(\b7_nYJ_BFM[301] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[302] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_286 (.A(b3_PLF_16_net_1), .B(
        b3_PLF_15_net_1), .C(b3_PLF_14_net_1), .D(b3_PLF_13_net_1), .Y(
        b3_PLF_286_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_129 (.A(\b7_nYJ_BFM[311] ), .B(
        \b7_nYJ_BFM[184] ), .C(\b7_vFW_PlM[310] ), .D(
        \b7_vFW_PlM[183] ), .Y(b3_PLF_129_net_1));
    SLE \genblk9.b7_nYJ_BFM[74]  (.D(\b7_nYJ_BFM[73] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[74] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_140 (.A(\b7_nYJ_BFM[200] ), .B(
        \b7_nYJ_BFM[73] ), .C(\b7_vFW_PlM[199] ), .D(\b7_vFW_PlM[72] ), 
        .Y(b3_PLF_140_net_1));
    SLE \genblk9.b7_nYJ_BFM[356]  (.D(\b7_nYJ_BFM[355] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[356] ));
    SLE \genblk9.b7_nYJ_BFM[301]  (.D(\b7_nYJ_BFM[300] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[301] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_154 (.A(\b7_nYJ_BFM[341] ), .B(
        \b7_nYJ_BFM[85] ), .C(\b7_vFW_PlM[340] ), .D(\b7_vFW_PlM[84] ), 
        .Y(b3_PLF_154_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_79 (.A(\b7_nYJ_BFM[284] ), .B(
        \b7_nYJ_BFM[173] ), .C(\b7_vFW_PlM[283] ), .D(
        \b7_vFW_PlM[172] ), .Y(b3_PLF_79_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_143 (.A(\b7_nYJ_BFM[196] ), .B(
        \b7_nYJ_BFM[69] ), .C(\b7_vFW_PlM[195] ), .D(\b7_vFW_PlM[68] ), 
        .Y(b3_PLF_143_net_1));
    SLE \genblk9.b7_nYJ_BFM[207]  (.D(\b7_nYJ_BFM[206] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[207] ));
    SLE \genblk9.b7_nYJ_BFM[93]  (.D(\b7_nYJ_BFM[92] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[93] ));
    SLE \genblk9.b7_nYJ_BFM[127]  (.D(\b7_nYJ_BFM[126] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[127] ));
    SLE \b12_PSyi_KyDbLbb[3]  (.D(\b12_2_St6KCa_jHv[3]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_184 (.A(\b7_nYJ_BFM[283] ), .B(
        \b7_nYJ_BFM[172] ), .C(\b7_vFW_PlM[282] ), .D(
        \b7_vFW_PlM[171] ), .Y(b3_PLF_184_net_1));
    SLE \genblk9.b7_nYJ_BFM[64]  (.D(\b7_nYJ_BFM[63] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[64] ));
    SLE \genblk9.b7_nYJ_BFM[250]  (.D(\b7_nYJ_BFM[249] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[250] ));
    CFG4 #( .INIT(16'h8000) )  b8_jAA_KlCO_0_sqmuxa (.A(
        \b12_2_St6KCa_jHv[3]_net_1 ), .B(\b12_2_St6KCa_jHv[4]_net_1 ), 
        .C(b8_jAA_KlCO_0_sqmuxa_8_net_1), .D(
        b8_jAA_KlCO_0_sqmuxa_4_net_1), .Y(b8_jAA_KlCO_0_sqmuxa_net_1));
    SLE \genblk9.b7_nYJ_BFM[263]  (.D(\b7_nYJ_BFM[262] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[263] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_92 (.A(\b7_nYJ_BFM[44] ), .B(
        \b7_nYJ_BFM[27] ), .C(\b7_vFW_PlM[43] ), .D(\b7_vFW_PlM[26] ), 
        .Y(b3_PLF_92_net_1));
    SLE \genblk9.b7_nYJ_BFM[243]  (.D(\b7_nYJ_BFM[242] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[243] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_326 (.A(b3_PLF_176_net_1), .B(
        b3_PLF_175_net_1), .C(b3_PLF_174_net_1), .D(b3_PLF_173_net_1), 
        .Y(b3_PLF_326_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_11 (.A(\b7_nYJ_BFM[151] ), .B(
        \b7_nYJ_BFM[24] ), .C(\b7_vFW_PlM[150] ), .D(\b7_vFW_PlM[23] ), 
        .Y(b3_PLF_11_net_1));
    SLE \genblk9.b7_nYJ_BFM[177]  (.D(\b7_nYJ_BFM[176] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[177] ));
    SLE \genblk9.b7_nYJ_BFM[327]  (.D(\b7_nYJ_BFM[326] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[327] ));
    SLE \genblk9.b7_nYJ_BFM[16]  (.D(\b7_nYJ_BFM[15] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[16] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_107 (.A(\b7_nYJ_BFM[150] ), .B(
        \b7_nYJ_BFM[23] ), .C(\b7_vFW_PlM[149] ), .D(\b7_vFW_PlM[22] ), 
        .Y(b3_PLF_107_net_1));
    SLE \genblk9.b7_nYJ_BFM[58]  (.D(\b7_nYJ_BFM[57] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[58] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_9 (.A(\b7_nYJ_BFM[282] ), .B(
        \b7_nYJ_BFM[26] ), .C(\b7_vFW_PlM[281] ), .D(\b7_vFW_PlM[25] ), 
        .Y(b3_PLF_9_net_1));
    SLE \genblk9.b7_nYJ_BFM[162]  (.D(\b7_nYJ_BFM[161] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[162] ));
    SLE \genblk9.b9_v_mzCDYXs[8]  (.D(b9_v_mzCDYXs_4), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[8] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNINN0G5[2]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[2] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_1), .S(\b9_v_mzCDYXs_RNINN0G5_S[2] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_2));
    SLE \genblk9.b7_nYJ_BFM[142]  (.D(\b7_nYJ_BFM[141] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[142] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_51 (.A(\b7_nYJ_BFM[322] ), .B(
        \b7_nYJ_BFM[66] ), .C(\b7_vFW_PlM[321] ), .D(\b7_vFW_PlM[65] ), 
        .Y(b3_PLF_51_net_1));
    SLE \genblk9.b7_nYJ_BFM[354]  (.D(\b7_nYJ_BFM[353] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[354] ));
    SLE \genblk9.b7_nYJ_BFM[328]  (.D(\b7_nYJ_BFM[327] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[328] ));
    SLE \genblk9.b7_nYJ_BFM[196]  (.D(\b7_nYJ_BFM[195] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[196] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_85 (.A(\b7_nYJ_BFM[372] ), .B(
        \b7_nYJ_BFM[245] ), .C(\b7_vFW_PlM[371] ), .D(
        \b7_vFW_PlM[244] ), .Y(b3_PLF_85_net_1));
    SLE \genblk9.b7_nYJ_BFM[20]  (.D(\b7_nYJ_BFM[19] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[20] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_299 (.A(b3_PLF_68_net_1), .B(
        b3_PLF_67_net_1), .C(b3_PLF_66_net_1), .D(b3_PLF_65_net_1), .Y(
        b3_PLF_299_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_65 (.A(\b7_nYJ_BFM[191] ), .B(
        \b7_nYJ_BFM[80] ), .C(\b7_vFW_PlM[190] ), .D(\b7_vFW_PlM[79] ), 
        .Y(b3_PLF_65_net_1));
    SLE \genblk9.b7_nYJ_BFM[38]  (.D(\b7_nYJ_BFM[37] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[38] ));
    SLE \genblk9.b7_nYJ_BFM[100]  (.D(\b7_nYJ_BFM[99] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[100] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIUDLP4[0]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[0] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_0_cy), .S(\b9_v_mzCDYXs_RNIUDLP4_S[0] )
        , .Y(), .FCO(b9_v_mzCDYXs_cry_0));
    SLE \genblk9.b7_nYJ_BFM[377]  (.D(\b7_nYJ_BFM[376] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[377] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_88 (.A(\b7_nYJ_BFM[368] ), .B(
        \b7_nYJ_BFM[241] ), .C(\b7_vFW_PlM[367] ), .D(
        \b7_vFW_PlM[240] ), .Y(b3_PLF_88_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_68 (.A(\b7_nYJ_BFM[251] ), .B(
        \b7_nYJ_BFM[12] ), .C(\b7_vFW_PlM[250] ), .D(\b7_vFW_PlM[11] ), 
        .Y(b3_PLF_68_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_30 (.A(\b7_nYJ_BFM[365] ), .B(
        \b7_nYJ_BFM[254] ), .C(\b7_vFW_PlM[364] ), .D(
        \b7_vFW_PlM[253] ), .Y(b3_PLF_30_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_102 (.A(\b7_nYJ_BFM[205] ), .B(
        \b7_nYJ_BFM[94] ), .C(\b7_vFW_PlM[204] ), .D(\b7_vFW_PlM[93] ), 
        .Y(b3_PLF_102_net_1));
    SLE \genblk9.b7_nYJ_BFM[94]  (.D(\b7_nYJ_BFM[93] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[94] ));
    SLE \genblk9.b7_nYJ_BFM[378]  (.D(\b7_nYJ_BFM[377] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[378] ));
    SLE \genblk9.b7_nYJ_BFM[117]  (.D(\b7_nYJ_BFM[116] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[117] ));
    SLE b8_jAA_KlCO (.D(VCC_net_1), .CLK(BW_clk_c), .EN(
        b8_jAA_KlCO_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b8_jAA_KlCO_net_1));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b9_v_mzCDYXs_RNIJKMC1[0]  (.A(
        \b9_v_mzCDYXs[4] ), .B(\b9_v_mzCDYXs[2] ), .C(
        \b9_v_mzCDYXs[1] ), .D(\b9_v_mzCDYXs[0] ), .Y(m9_e_5));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_137 (.A(\b7_nYJ_BFM[253] ), .B(
        \b7_nYJ_BFM[13] ), .C(\b7_vFW_PlM[252] ), .D(\b7_vFW_PlM[12] ), 
        .Y(b3_PLF_137_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_46 (.A(\b7_nYJ_BFM[328] ), .B(
        \b7_nYJ_BFM[201] ), .C(\b7_vFW_PlM[327] ), .D(
        \b7_vFW_PlM[200] ), .Y(b3_PLF_46_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[3]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNI5E6R5_S[3] ), .Y(b9_v_mzCDYXs));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_364 (.A(b3_PLF_328_net_1), .B(
        b3_PLF_327_net_1), .C(b3_PLF_326_net_1), .D(b3_PLF_325_net_1), 
        .Y(b3_PLF_364_net_1));
    b13_vFW_xNywD_EdR_383s_10s_1024s_0s_x_0 b3_SoW (.IICE_comm2iice({
        IICE_comm2iice_11}), .b12_2_St6KCa_jHv({
        \b12_2_St6KCa_jHv[9]_net_1 , \b12_2_St6KCa_jHv[8]_net_1 , 
        \b12_2_St6KCa_jHv[7]_net_1 , \b12_2_St6KCa_jHv[6]_net_1 , 
        \b12_2_St6KCa_jHv[5]_net_1 , \b12_2_St6KCa_jHv[4]_net_1 , 
        \b12_2_St6KCa_jHv[3]_net_1 , \b12_2_St6KCa_jHv[2]_net_1 , 
        \b12_2_St6KCa_jHv[1]_net_1 , \b12_2_St6KCa_jHv[0]_net_1 }), 
        .b7_vFW_PlM({\b7_vFW_PlM[376] , \b7_vFW_PlM[375] , 
        \b7_vFW_PlM[374] , \b7_vFW_PlM[373] , \b7_vFW_PlM[372] , 
        \b7_vFW_PlM[371] , \b7_vFW_PlM[370] , \b7_vFW_PlM[369] , 
        \b7_vFW_PlM[368] , \b7_vFW_PlM[367] , \b7_vFW_PlM[366] , 
        \b7_vFW_PlM[365] , \b7_vFW_PlM[364] , \b7_vFW_PlM[363] , 
        \b7_vFW_PlM[362] , \b7_vFW_PlM[361] , \b7_vFW_PlM[360] , 
        \b7_vFW_PlM[359] , \b7_vFW_PlM[358] , \b7_vFW_PlM[357] , 
        \b7_vFW_PlM[356] , \b7_vFW_PlM[355] , \b7_vFW_PlM[354] , 
        \b7_vFW_PlM[353] , \b7_vFW_PlM[352] , \b7_vFW_PlM[351] , 
        \b7_vFW_PlM[350] , \b7_vFW_PlM[349] , \b7_vFW_PlM[348] , 
        \b7_vFW_PlM[347] , \b7_vFW_PlM[346] , \b7_vFW_PlM[345] , 
        \b7_vFW_PlM[344] , \b7_vFW_PlM[343] , \b7_vFW_PlM[342] , 
        \b7_vFW_PlM[341] , \b7_vFW_PlM[340] , \b7_vFW_PlM[339] , 
        \b7_vFW_PlM[338] , \b7_vFW_PlM[337] , \b7_vFW_PlM[336] , 
        \b7_vFW_PlM[335] , \b7_vFW_PlM[334] , \b7_vFW_PlM[333] , 
        \b7_vFW_PlM[332] , \b7_vFW_PlM[331] , \b7_vFW_PlM[330] , 
        \b7_vFW_PlM[329] , \b7_vFW_PlM[328] , \b7_vFW_PlM[327] , 
        \b7_vFW_PlM[326] , \b7_vFW_PlM[325] , \b7_vFW_PlM[324] , 
        \b7_vFW_PlM[323] , \b7_vFW_PlM[322] , \b7_vFW_PlM[321] , 
        \b7_vFW_PlM[320] , \b7_vFW_PlM[319] , \b7_vFW_PlM[318] , 
        \b7_vFW_PlM[317] , \b7_vFW_PlM[316] , \b7_vFW_PlM[315] , 
        \b7_vFW_PlM[314] , \b7_vFW_PlM[313] , \b7_vFW_PlM[312] , 
        \b7_vFW_PlM[311] , \b7_vFW_PlM[310] , \b7_vFW_PlM[309] , 
        \b7_vFW_PlM[308] , \b7_vFW_PlM[307] , \b7_vFW_PlM[306] , 
        \b7_vFW_PlM[305] , \b7_vFW_PlM[304] , \b7_vFW_PlM[303] , 
        \b7_vFW_PlM[302] , \b7_vFW_PlM[301] , \b7_vFW_PlM[300] , 
        \b7_vFW_PlM[299] , \b7_vFW_PlM[298] , \b7_vFW_PlM[297] , 
        \b7_vFW_PlM[296] , \b7_vFW_PlM[295] , \b7_vFW_PlM[294] , 
        \b7_vFW_PlM[293] , \b7_vFW_PlM[292] , \b7_vFW_PlM[291] , 
        \b7_vFW_PlM[290] , \b7_vFW_PlM[289] , \b7_vFW_PlM[288] , 
        \b7_vFW_PlM[287] , \b7_vFW_PlM[286] , \b7_vFW_PlM[285] , 
        \b7_vFW_PlM[284] , \b7_vFW_PlM[283] , \b7_vFW_PlM[282] , 
        \b7_vFW_PlM[281] , \b7_vFW_PlM[280] , \b7_vFW_PlM[279] , 
        \b7_vFW_PlM[278] , \b7_vFW_PlM[277] , \b7_vFW_PlM[276] , 
        \b7_vFW_PlM[275] , \b7_vFW_PlM[274] , \b7_vFW_PlM[273] , 
        \b7_vFW_PlM[272] , \b7_vFW_PlM[271] , \b7_vFW_PlM[270] , 
        \b7_vFW_PlM[269] , \b7_vFW_PlM[268] , \b7_vFW_PlM[267] , 
        \b7_vFW_PlM[266] , \b7_vFW_PlM[265] , \b7_vFW_PlM[264] , 
        \b7_vFW_PlM[263] , \b7_vFW_PlM[262] , \b7_vFW_PlM[261] , 
        \b7_vFW_PlM[260] , \b7_vFW_PlM[259] , \b7_vFW_PlM[258] , 
        \b7_vFW_PlM[257] , \b7_vFW_PlM[256] , \b7_vFW_PlM[255] , 
        \b7_vFW_PlM[254] , \b7_vFW_PlM[253] , \b7_vFW_PlM[252] , 
        \b7_vFW_PlM[251] , \b7_vFW_PlM[250] , \b7_vFW_PlM[249] , 
        \b7_vFW_PlM[248] , \b7_vFW_PlM[247] , \b7_vFW_PlM[246] , 
        \b7_vFW_PlM[245] , \b7_vFW_PlM[244] , \b7_vFW_PlM[243] , 
        \b7_vFW_PlM[242] , \b7_vFW_PlM[241] , \b7_vFW_PlM[240] , 
        \b7_vFW_PlM[239] , \b7_vFW_PlM[238] , \b7_vFW_PlM[237] , 
        \b7_vFW_PlM[236] , \b7_vFW_PlM[235] , \b7_vFW_PlM[234] , 
        \b7_vFW_PlM[233] , \b7_vFW_PlM[232] , \b7_vFW_PlM[231] , 
        \b7_vFW_PlM[230] , \b7_vFW_PlM[229] , \b7_vFW_PlM[228] , 
        \b7_vFW_PlM[227] , \b7_vFW_PlM[226] , \b7_vFW_PlM[225] , 
        \b7_vFW_PlM[224] , \b7_vFW_PlM[223] , \b7_vFW_PlM[222] , 
        \b7_vFW_PlM[221] , \b7_vFW_PlM[220] , \b7_vFW_PlM[219] , 
        \b7_vFW_PlM[218] , \b7_vFW_PlM[217] , \b7_vFW_PlM[216] , 
        \b7_vFW_PlM[215] , \b7_vFW_PlM[214] , \b7_vFW_PlM[213] , 
        \b7_vFW_PlM[212] , \b7_vFW_PlM[211] , \b7_vFW_PlM[210] , 
        \b7_vFW_PlM[209] , \b7_vFW_PlM[208] , \b7_vFW_PlM[207] , 
        \b7_vFW_PlM[206] , \b7_vFW_PlM[205] , \b7_vFW_PlM[204] , 
        \b7_vFW_PlM[203] , \b7_vFW_PlM[202] , \b7_vFW_PlM[201] , 
        \b7_vFW_PlM[200] , \b7_vFW_PlM[199] , \b7_vFW_PlM[198] , 
        \b7_vFW_PlM[197] , \b7_vFW_PlM[196] , \b7_vFW_PlM[195] , 
        \b7_vFW_PlM[194] , \b7_vFW_PlM[193] , \b7_vFW_PlM[192] , 
        \b7_vFW_PlM[191] , \b7_vFW_PlM[190] , \b7_vFW_PlM[189] , 
        \b7_vFW_PlM[188] , \b7_vFW_PlM[187] , \b7_vFW_PlM[186] , 
        \b7_vFW_PlM[185] , \b7_vFW_PlM[184] , \b7_vFW_PlM[183] , 
        \b7_vFW_PlM[182] , \b7_vFW_PlM[181] , \b7_vFW_PlM[180] , 
        \b7_vFW_PlM[179] , \b7_vFW_PlM[178] , \b7_vFW_PlM[177] , 
        \b7_vFW_PlM[176] , \b7_vFW_PlM[175] , \b7_vFW_PlM[174] , 
        \b7_vFW_PlM[173] , \b7_vFW_PlM[172] , \b7_vFW_PlM[171] , 
        \b7_vFW_PlM[170] , \b7_vFW_PlM[169] , \b7_vFW_PlM[168] , 
        \b7_vFW_PlM[167] , \b7_vFW_PlM[166] , \b7_vFW_PlM[165] , 
        \b7_vFW_PlM[164] , \b7_vFW_PlM[163] , \b7_vFW_PlM[162] , 
        \b7_vFW_PlM[161] , \b7_vFW_PlM[160] , \b7_vFW_PlM[159] , 
        \b7_vFW_PlM[158] , \b7_vFW_PlM[157] , \b7_vFW_PlM[156] , 
        \b7_vFW_PlM[155] , \b7_vFW_PlM[154] , \b7_vFW_PlM[153] , 
        \b7_vFW_PlM[152] , \b7_vFW_PlM[151] , \b7_vFW_PlM[150] , 
        \b7_vFW_PlM[149] , \b7_vFW_PlM[148] , \b7_vFW_PlM[147] , 
        \b7_vFW_PlM[146] , \b7_vFW_PlM[145] , \b7_vFW_PlM[144] , 
        \b7_vFW_PlM[143] , \b7_vFW_PlM[142] , \b7_vFW_PlM[141] , 
        \b7_vFW_PlM[140] , \b7_vFW_PlM[139] , \b7_vFW_PlM[138] , 
        \b7_vFW_PlM[137] , \b7_vFW_PlM[136] , \b7_vFW_PlM[135] , 
        \b7_vFW_PlM[134] , \b7_vFW_PlM[133] , \b7_vFW_PlM[132] , 
        \b7_vFW_PlM[131] , \b7_vFW_PlM[130] , \b7_vFW_PlM[129] , 
        \b7_vFW_PlM[128] , \b7_vFW_PlM[127] , \b7_vFW_PlM[126] , 
        \b7_vFW_PlM[125] , \b7_vFW_PlM[124] , \b7_vFW_PlM[123] , 
        \b7_vFW_PlM[122] , \b7_vFW_PlM[121] , \b7_vFW_PlM[120] , 
        \b7_vFW_PlM[119] , \b7_vFW_PlM[118] , \b7_vFW_PlM[117] , 
        \b7_vFW_PlM[116] , \b7_vFW_PlM[115] , \b7_vFW_PlM[114] , 
        \b7_vFW_PlM[113] , \b7_vFW_PlM[112] , \b7_vFW_PlM[111] , 
        \b7_vFW_PlM[110] , \b7_vFW_PlM[109] , \b7_vFW_PlM[108] , 
        \b7_vFW_PlM[107] , \b7_vFW_PlM[106] , \b7_vFW_PlM[105] , 
        \b7_vFW_PlM[104] , \b7_vFW_PlM[103] , \b7_vFW_PlM[102] , 
        \b7_vFW_PlM[101] , \b7_vFW_PlM[100] , \b7_vFW_PlM[99] , 
        \b7_vFW_PlM[98] , \b7_vFW_PlM[97] , \b7_vFW_PlM[96] , 
        \b7_vFW_PlM[95] , \b7_vFW_PlM[94] , \b7_vFW_PlM[93] , 
        \b7_vFW_PlM[92] , \b7_vFW_PlM[91] , \b7_vFW_PlM[90] , 
        \b7_vFW_PlM[89] , \b7_vFW_PlM[88] , \b7_vFW_PlM[87] , 
        \b7_vFW_PlM[86] , \b7_vFW_PlM[85] , \b7_vFW_PlM[84] , 
        \b7_vFW_PlM[83] , \b7_vFW_PlM[82] , \b7_vFW_PlM[81] , 
        \b7_vFW_PlM[80] , \b7_vFW_PlM[79] , \b7_vFW_PlM[78] , 
        \b7_vFW_PlM[77] , \b7_vFW_PlM[76] , \b7_vFW_PlM[75] , 
        \b7_vFW_PlM[74] , \b7_vFW_PlM[73] , \b7_vFW_PlM[72] , 
        \b7_vFW_PlM[71] , \b7_vFW_PlM[70] , \b7_vFW_PlM[69] , 
        \b7_vFW_PlM[68] , \b7_vFW_PlM[67] , \b7_vFW_PlM[66] , 
        \b7_vFW_PlM[65] , \b7_vFW_PlM[64] , \b7_vFW_PlM[63] , 
        \b7_vFW_PlM[62] , \b7_vFW_PlM[61] , \b7_vFW_PlM[60] , 
        \b7_vFW_PlM[59] , \b7_vFW_PlM[58] , \b7_vFW_PlM[57] , 
        \b7_vFW_PlM[56] , \b7_vFW_PlM[55] , \b7_vFW_PlM[54] , 
        \b7_vFW_PlM[53] , \b7_vFW_PlM[52] , \b7_vFW_PlM[51] , 
        \b7_vFW_PlM[50] , \b7_vFW_PlM[49] , \b7_vFW_PlM[48] , 
        \b7_vFW_PlM[47] , \b7_vFW_PlM[46] , \b7_vFW_PlM[45] , 
        \b7_vFW_PlM[44] , \b7_vFW_PlM[43] , \b7_vFW_PlM[42] , 
        \b7_vFW_PlM[41] , \b7_vFW_PlM[40] , \b7_vFW_PlM[39] , 
        \b7_vFW_PlM[38] , \b7_vFW_PlM[37] , \b7_vFW_PlM[36] , 
        \b7_vFW_PlM[35] , \b7_vFW_PlM[34] , \b7_vFW_PlM[33] , 
        \b7_vFW_PlM[32] , \b7_vFW_PlM[31] , \b7_vFW_PlM[30] , 
        \b7_vFW_PlM[29] , \b7_vFW_PlM[28] , \b7_vFW_PlM[27] , 
        \b7_vFW_PlM[26] , \b7_vFW_PlM[25] , \b7_vFW_PlM[24] , 
        \b7_vFW_PlM[23] , \b7_vFW_PlM[22] , \b7_vFW_PlM[21] , 
        \b7_vFW_PlM[20] , \b7_vFW_PlM[19] , \b7_vFW_PlM[18] , 
        \b7_vFW_PlM[17] , \b7_vFW_PlM[16] , \b7_vFW_PlM[15] , 
        \b7_vFW_PlM[14] , \b7_vFW_PlM[13] , \b7_vFW_PlM[12] , 
        \b7_vFW_PlM[11] , \b7_vFW_PlM[10] , \b7_vFW_PlM[9] , 
        \b7_vFW_PlM[8] , \b7_vFW_PlM[7] , \b7_vFW_PlM[6] , 
        \b7_vFW_PlM[5] , \b7_vFW_PlM[4] , \b7_vFW_PlM[3] , 
        \b7_vFW_PlM[2] , \b7_vFW_PlM[1] , \b7_vFW_PlM[0] }), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[376], b11_OFWNT9L_8tZ[375], 
        b11_OFWNT9L_8tZ[374], b11_OFWNT9L_8tZ[373], 
        b11_OFWNT9L_8tZ[372], b11_OFWNT9L_8tZ[371], 
        b11_OFWNT9L_8tZ[370], b11_OFWNT9L_8tZ[369], 
        b11_OFWNT9L_8tZ[368], b11_OFWNT9L_8tZ[367], 
        b11_OFWNT9L_8tZ[366], b11_OFWNT9L_8tZ[365], 
        b11_OFWNT9L_8tZ[364], b11_OFWNT9L_8tZ[363], 
        b11_OFWNT9L_8tZ[362], b11_OFWNT9L_8tZ[361], 
        b11_OFWNT9L_8tZ[360], b11_OFWNT9L_8tZ[359], 
        b11_OFWNT9L_8tZ[358], b11_OFWNT9L_8tZ[357], 
        b11_OFWNT9L_8tZ[356], b11_OFWNT9L_8tZ[355], 
        b11_OFWNT9L_8tZ[354], b11_OFWNT9L_8tZ[353], 
        b11_OFWNT9L_8tZ[352], b11_OFWNT9L_8tZ[351], 
        b11_OFWNT9L_8tZ[350], b11_OFWNT9L_8tZ[349], 
        b11_OFWNT9L_8tZ[348], b11_OFWNT9L_8tZ[347], 
        b11_OFWNT9L_8tZ[346], b11_OFWNT9L_8tZ[345], 
        b11_OFWNT9L_8tZ[344], b11_OFWNT9L_8tZ[343], 
        b11_OFWNT9L_8tZ[342], b11_OFWNT9L_8tZ[341], 
        b11_OFWNT9L_8tZ[340], b11_OFWNT9L_8tZ[339], 
        b11_OFWNT9L_8tZ[338], b11_OFWNT9L_8tZ[337], 
        b11_OFWNT9L_8tZ[336], b11_OFWNT9L_8tZ[335], 
        b11_OFWNT9L_8tZ[334], b11_OFWNT9L_8tZ[333], 
        b11_OFWNT9L_8tZ[332], b11_OFWNT9L_8tZ[331], 
        b11_OFWNT9L_8tZ[330], b11_OFWNT9L_8tZ[329], 
        b11_OFWNT9L_8tZ[328], b11_OFWNT9L_8tZ[327], 
        b11_OFWNT9L_8tZ[326], b11_OFWNT9L_8tZ[325], 
        b11_OFWNT9L_8tZ[324], b11_OFWNT9L_8tZ[323], 
        b11_OFWNT9L_8tZ[322], b11_OFWNT9L_8tZ[321], 
        b11_OFWNT9L_8tZ[320], b11_OFWNT9L_8tZ[319], 
        b11_OFWNT9L_8tZ[318], b11_OFWNT9L_8tZ[317], 
        b11_OFWNT9L_8tZ[316], b11_OFWNT9L_8tZ[315], 
        b11_OFWNT9L_8tZ[314], b11_OFWNT9L_8tZ[313], 
        b11_OFWNT9L_8tZ[312], b11_OFWNT9L_8tZ[311], 
        b11_OFWNT9L_8tZ[310], b11_OFWNT9L_8tZ[309], 
        b11_OFWNT9L_8tZ[308], b11_OFWNT9L_8tZ[307], 
        b11_OFWNT9L_8tZ[306], b11_OFWNT9L_8tZ[305], 
        b11_OFWNT9L_8tZ[304], b11_OFWNT9L_8tZ[303], 
        b11_OFWNT9L_8tZ[302], b11_OFWNT9L_8tZ[301], 
        b11_OFWNT9L_8tZ[300], b11_OFWNT9L_8tZ[299], 
        b11_OFWNT9L_8tZ[298], b11_OFWNT9L_8tZ[297], 
        b11_OFWNT9L_8tZ[296], b11_OFWNT9L_8tZ[295], 
        b11_OFWNT9L_8tZ[294], b11_OFWNT9L_8tZ[293], 
        b11_OFWNT9L_8tZ[292], b11_OFWNT9L_8tZ[291], 
        b11_OFWNT9L_8tZ[290], b11_OFWNT9L_8tZ[289], 
        b11_OFWNT9L_8tZ[288], b11_OFWNT9L_8tZ[287], 
        b11_OFWNT9L_8tZ[286], b11_OFWNT9L_8tZ[285], 
        b11_OFWNT9L_8tZ[284], b11_OFWNT9L_8tZ[283], 
        b11_OFWNT9L_8tZ[282], b11_OFWNT9L_8tZ[281], 
        b11_OFWNT9L_8tZ[280], b11_OFWNT9L_8tZ[279], 
        b11_OFWNT9L_8tZ[278], b11_OFWNT9L_8tZ[277], 
        b11_OFWNT9L_8tZ[276], b11_OFWNT9L_8tZ[275], 
        b11_OFWNT9L_8tZ[274], b11_OFWNT9L_8tZ[273], 
        b11_OFWNT9L_8tZ[272], b11_OFWNT9L_8tZ[271], 
        b11_OFWNT9L_8tZ[270], b11_OFWNT9L_8tZ[269], 
        b11_OFWNT9L_8tZ[268], b11_OFWNT9L_8tZ[267], 
        b11_OFWNT9L_8tZ[266], b11_OFWNT9L_8tZ[265], 
        b11_OFWNT9L_8tZ[264], b11_OFWNT9L_8tZ[263], 
        b11_OFWNT9L_8tZ[262], b11_OFWNT9L_8tZ[261], 
        b11_OFWNT9L_8tZ[260], b11_OFWNT9L_8tZ[259], 
        b11_OFWNT9L_8tZ[258], b11_OFWNT9L_8tZ[257], 
        b11_OFWNT9L_8tZ[256], b11_OFWNT9L_8tZ[255], 
        b11_OFWNT9L_8tZ[254], b11_OFWNT9L_8tZ[253], 
        b11_OFWNT9L_8tZ[252], b11_OFWNT9L_8tZ[251], 
        b11_OFWNT9L_8tZ[250], b11_OFWNT9L_8tZ[249], 
        b11_OFWNT9L_8tZ[248], b11_OFWNT9L_8tZ[247], 
        b11_OFWNT9L_8tZ[246], b11_OFWNT9L_8tZ[245], 
        b11_OFWNT9L_8tZ[244], b11_OFWNT9L_8tZ[243], 
        b11_OFWNT9L_8tZ[242], b11_OFWNT9L_8tZ[241], 
        b11_OFWNT9L_8tZ[240], b11_OFWNT9L_8tZ[239], 
        b11_OFWNT9L_8tZ[238], b11_OFWNT9L_8tZ[237], 
        b11_OFWNT9L_8tZ[236], b11_OFWNT9L_8tZ[235], 
        b11_OFWNT9L_8tZ[234], b11_OFWNT9L_8tZ[233], 
        b11_OFWNT9L_8tZ[232], b11_OFWNT9L_8tZ[231], 
        b11_OFWNT9L_8tZ[230], b11_OFWNT9L_8tZ[229], 
        b11_OFWNT9L_8tZ[228], b11_OFWNT9L_8tZ[227], 
        b11_OFWNT9L_8tZ[226], b11_OFWNT9L_8tZ[225], 
        b11_OFWNT9L_8tZ[224], b11_OFWNT9L_8tZ[223], 
        b11_OFWNT9L_8tZ[222], b11_OFWNT9L_8tZ[221], 
        b11_OFWNT9L_8tZ[220], b11_OFWNT9L_8tZ[219], 
        b11_OFWNT9L_8tZ[218], b11_OFWNT9L_8tZ[217], 
        b11_OFWNT9L_8tZ[216], b11_OFWNT9L_8tZ[215], 
        b11_OFWNT9L_8tZ[214], b11_OFWNT9L_8tZ[213], 
        b11_OFWNT9L_8tZ[212], b11_OFWNT9L_8tZ[211], 
        b11_OFWNT9L_8tZ[210], b11_OFWNT9L_8tZ[209], 
        b11_OFWNT9L_8tZ[208], b11_OFWNT9L_8tZ[207], 
        b11_OFWNT9L_8tZ[206], b11_OFWNT9L_8tZ[205], 
        b11_OFWNT9L_8tZ[204], b11_OFWNT9L_8tZ[203], 
        b11_OFWNT9L_8tZ[202], b11_OFWNT9L_8tZ[201], 
        b11_OFWNT9L_8tZ[200], b11_OFWNT9L_8tZ[199], 
        b11_OFWNT9L_8tZ[198], b11_OFWNT9L_8tZ[197], 
        b11_OFWNT9L_8tZ[196], b11_OFWNT9L_8tZ[195], 
        b11_OFWNT9L_8tZ[194], b11_OFWNT9L_8tZ[193], 
        b11_OFWNT9L_8tZ[192], b11_OFWNT9L_8tZ[191], 
        b11_OFWNT9L_8tZ[190], b11_OFWNT9L_8tZ[189], 
        b11_OFWNT9L_8tZ[188], b11_OFWNT9L_8tZ[187], 
        b11_OFWNT9L_8tZ[186], b11_OFWNT9L_8tZ[185], 
        b11_OFWNT9L_8tZ[184], b11_OFWNT9L_8tZ[183], 
        b11_OFWNT9L_8tZ[182], b11_OFWNT9L_8tZ[181], 
        b11_OFWNT9L_8tZ[180], b11_OFWNT9L_8tZ[179], 
        b11_OFWNT9L_8tZ[178], b11_OFWNT9L_8tZ[177], 
        b11_OFWNT9L_8tZ[176], b11_OFWNT9L_8tZ[175], 
        b11_OFWNT9L_8tZ[174], b11_OFWNT9L_8tZ[173], 
        b11_OFWNT9L_8tZ[172], b11_OFWNT9L_8tZ[171], 
        b11_OFWNT9L_8tZ[170], b11_OFWNT9L_8tZ[169], 
        b11_OFWNT9L_8tZ[168], b11_OFWNT9L_8tZ[167], 
        b11_OFWNT9L_8tZ[166], b11_OFWNT9L_8tZ[165], 
        b11_OFWNT9L_8tZ[164], b11_OFWNT9L_8tZ[163], 
        b11_OFWNT9L_8tZ[162], b11_OFWNT9L_8tZ[161], 
        b11_OFWNT9L_8tZ[160], b11_OFWNT9L_8tZ[159], 
        b11_OFWNT9L_8tZ[158], b11_OFWNT9L_8tZ[157], 
        b11_OFWNT9L_8tZ[156], b11_OFWNT9L_8tZ[155], 
        b11_OFWNT9L_8tZ[154], b11_OFWNT9L_8tZ[153], 
        b11_OFWNT9L_8tZ[152], b11_OFWNT9L_8tZ[151], 
        b11_OFWNT9L_8tZ[150], b11_OFWNT9L_8tZ[149], 
        b11_OFWNT9L_8tZ[148], b11_OFWNT9L_8tZ[147], 
        b11_OFWNT9L_8tZ[146], b11_OFWNT9L_8tZ[145], 
        b11_OFWNT9L_8tZ[144], b11_OFWNT9L_8tZ[143], 
        b11_OFWNT9L_8tZ[142], b11_OFWNT9L_8tZ[141], 
        b11_OFWNT9L_8tZ[140], b11_OFWNT9L_8tZ[139], 
        b11_OFWNT9L_8tZ[138], b11_OFWNT9L_8tZ[137], 
        b11_OFWNT9L_8tZ[136], b11_OFWNT9L_8tZ[135], 
        b11_OFWNT9L_8tZ[134], b11_OFWNT9L_8tZ[133], 
        b11_OFWNT9L_8tZ[132], b11_OFWNT9L_8tZ[131], 
        b11_OFWNT9L_8tZ[130], b11_OFWNT9L_8tZ[129], 
        b11_OFWNT9L_8tZ[128], b11_OFWNT9L_8tZ[127], 
        b11_OFWNT9L_8tZ[126], b11_OFWNT9L_8tZ[125], 
        b11_OFWNT9L_8tZ[124], b11_OFWNT9L_8tZ[123], 
        b11_OFWNT9L_8tZ[122], b11_OFWNT9L_8tZ[121], 
        b11_OFWNT9L_8tZ[120], b11_OFWNT9L_8tZ[119], 
        b11_OFWNT9L_8tZ[118], b11_OFWNT9L_8tZ[117], 
        b11_OFWNT9L_8tZ[116], b11_OFWNT9L_8tZ[115], 
        b11_OFWNT9L_8tZ[114], b11_OFWNT9L_8tZ[113], 
        b11_OFWNT9L_8tZ[112], b11_OFWNT9L_8tZ[111], 
        b11_OFWNT9L_8tZ[110], b11_OFWNT9L_8tZ[109], 
        b11_OFWNT9L_8tZ[108], b11_OFWNT9L_8tZ[107], 
        b11_OFWNT9L_8tZ[106], b11_OFWNT9L_8tZ[105], 
        b11_OFWNT9L_8tZ[104], b11_OFWNT9L_8tZ[103], 
        b11_OFWNT9L_8tZ[102], b11_OFWNT9L_8tZ[101], 
        b11_OFWNT9L_8tZ[100], b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], 
        b11_OFWNT9L_8tZ[97], b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], 
        b11_OFWNT9L_8tZ[94], b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], 
        b11_OFWNT9L_8tZ[91], b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], 
        b11_OFWNT9L_8tZ[88], b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], 
        b11_OFWNT9L_8tZ[85], b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], 
        b11_OFWNT9L_8tZ[82], b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], 
        b11_OFWNT9L_8tZ[79], b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], 
        b11_OFWNT9L_8tZ[76], b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], 
        b11_OFWNT9L_8tZ[73], b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], 
        b11_OFWNT9L_8tZ[70], b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], 
        b11_OFWNT9L_8tZ[67], b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], 
        b11_OFWNT9L_8tZ[64], b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], 
        b11_OFWNT9L_8tZ[61], b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], 
        b11_OFWNT9L_8tZ[58], b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], 
        b11_OFWNT9L_8tZ[55], b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], 
        b11_OFWNT9L_8tZ[52], b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], 
        b11_OFWNT9L_8tZ[49], b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], 
        b11_OFWNT9L_8tZ[46], b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], 
        b11_OFWNT9L_8tZ[43], b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], 
        b11_OFWNT9L_8tZ[40], b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], 
        b11_OFWNT9L_8tZ[37], b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], 
        b11_OFWNT9L_8tZ[34], b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], 
        b11_OFWNT9L_8tZ[31], b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], 
        b11_OFWNT9L_8tZ[28], b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], 
        b11_OFWNT9L_8tZ[25], b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], 
        b11_OFWNT9L_8tZ[22], b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], 
        b11_OFWNT9L_8tZ[19], b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], 
        b11_OFWNT9L_8tZ[16], b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], 
        b11_OFWNT9L_8tZ[13], b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], 
        b11_OFWNT9L_8tZ[10], b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], 
        b11_OFWNT9L_8tZ[7], b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], 
        b11_OFWNT9L_8tZ[4], b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], 
        b11_OFWNT9L_8tZ[1], b11_OFWNT9L_8tZ[0]}), .b9_v_mzCDYXs_2(
        b9_v_mzCDYXs_2), .b9_v_mzCDYXs_1(b9_v_mzCDYXs_1), 
        .b9_v_mzCDYXs_0(b9_v_mzCDYXs_0), .b9_v_mzCDYXs(b9_v_mzCDYXs), 
        .b9_v_mzCDYXs_8(b9_v_mzCDYXs_8), .b9_v_mzCDYXs_7(
        b9_v_mzCDYXs_7), .b9_v_mzCDYXs_6(b9_v_mzCDYXs_6), 
        .b9_v_mzCDYXs_5(b9_v_mzCDYXs_5), .b9_v_mzCDYXs_4(
        b9_v_mzCDYXs_4), .b9_v_mzCDYXs_3(b9_v_mzCDYXs_3), .BW_clk_c(
        BW_clk_c), .b4_2o_z(b4_2o_z));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_17 (.A(\b7_nYJ_BFM[127] ), .B(
        \b7_nYJ_BFM[16] ), .C(\b7_vFW_PlM[126] ), .D(\b7_vFW_PlM[15] ), 
        .Y(b3_PLF_17_net_1));
    SLE \genblk9.b7_nYJ_BFM[317]  (.D(\b7_nYJ_BFM[316] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[317] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[4]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_4_S), .Y(b12_2_St6KCa_jHv_3));
    SLE \genblk9.b7_nYJ_BFM[45]  (.D(\b7_nYJ_BFM[44] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[45] ));
    SLE \genblk9.b7_nYJ_BFM[329]  (.D(\b7_nYJ_BFM[328] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[329] ));
    SLE \genblk9.b7_nYJ_BFM[318]  (.D(\b7_nYJ_BFM[317] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[318] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_57 (.A(\b7_nYJ_BFM[346] ), .B(
        \b7_nYJ_BFM[90] ), .C(\b7_vFW_PlM[345] ), .D(\b7_vFW_PlM[89] ), 
        .Y(b3_PLF_57_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_33 (.A(\b7_nYJ_BFM[314] ), .B(
        \b7_nYJ_BFM[58] ), .C(\b7_vFW_PlM[313] ), .D(\b7_vFW_PlM[57] ), 
        .Y(b3_PLF_33_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_132 (.A(\b7_nYJ_BFM[307] ), .B(
        \b7_nYJ_BFM[180] ), .C(\b7_vFW_PlM[306] ), .D(
        \b7_vFW_PlM[179] ), .Y(b3_PLF_132_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_22 (.A(\b7_nYJ_BFM[296] ), .B(
        \b7_nYJ_BFM[169] ), .C(\b7_vFW_PlM[295] ), .D(
        \b7_vFW_PlM[168] ), .Y(b3_PLF_22_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_362 (.A(b3_PLF_320_net_1), .B(
        b3_PLF_319_net_1), .C(b3_PLF_318_net_1), .D(b3_PLF_317_net_1), 
        .Y(b3_PLF_362_net_1));
    SLE \genblk9.b7_nYJ_BFM[225]  (.D(\b7_nYJ_BFM[224] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[225] ));
    b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0 virOut (.IICE_comm2iice_11(
        IICE_comm2iice_11), .IICE_comm2iice_9(IICE_comm2iice_9), 
        .IICE_comm2iice_1(IICE_comm2iice_1), .IICE_comm2iice_3(
        IICE_comm2iice_3), .IICE_comm2iice_2(IICE_comm2iice_2), 
        .IICE_comm2iice_4(IICE_comm2iice_4), .IICE_comm2iice_0(
        IICE_comm2iice_0), .IICE_comm2iice_5(IICE_comm2iice_5), 
        .IICE_comm2iice_6(IICE_comm2iice_6), .b4_ycsM(b4_ycsM), 
        .un1_b13_PLF_2grFt_FH911_i_a2_0_2(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .N_21(N_21), .un1_b5_OvyH3(
        un1_b5_OvyH3));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_2 (.A(\b7_nYJ_BFM[131] ), .B(
        \b7_nYJ_BFM[4] ), .C(\b7_vFW_PlM[130] ), .D(\b7_vFW_PlM[3] ), 
        .Y(b3_PLF_2_net_1));
    SLE \genblk9.b7_nYJ_BFM[187]  (.D(\b7_nYJ_BFM[186] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[187] ));
    SLE \genblk9.b7_nYJ_BFM[379]  (.D(\b7_nYJ_BFM[378] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[379] ));
    SLE \genblk9.b7_nYJ_BFM[352]  (.D(\b7_nYJ_BFM[351] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[352] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIK5C66[4]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[4] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_3), .S(\b9_v_mzCDYXs_RNIK5C66_S[4] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_4));
    b11_SoWyP0zEFKY_383s_0s_6s_0s_2s_2s_0s_0s_2s_0s_x_0 b6_SoWyQD (
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[376], b11_OFWNT9L_8tZ[375], 
        b11_OFWNT9L_8tZ[374], b11_OFWNT9L_8tZ[373], 
        b11_OFWNT9L_8tZ[372], b11_OFWNT9L_8tZ[371], 
        b11_OFWNT9L_8tZ[370], b11_OFWNT9L_8tZ[369], 
        b11_OFWNT9L_8tZ[368], b11_OFWNT9L_8tZ[367], 
        b11_OFWNT9L_8tZ[366], b11_OFWNT9L_8tZ[365], 
        b11_OFWNT9L_8tZ[364], b11_OFWNT9L_8tZ[363], 
        b11_OFWNT9L_8tZ[362], b11_OFWNT9L_8tZ[361], 
        b11_OFWNT9L_8tZ[360], b11_OFWNT9L_8tZ[359], 
        b11_OFWNT9L_8tZ[358], b11_OFWNT9L_8tZ[357], 
        b11_OFWNT9L_8tZ[356], b11_OFWNT9L_8tZ[355], 
        b11_OFWNT9L_8tZ[354], b11_OFWNT9L_8tZ[353], 
        b11_OFWNT9L_8tZ[352], b11_OFWNT9L_8tZ[351], 
        b11_OFWNT9L_8tZ[350], b11_OFWNT9L_8tZ[349], 
        b11_OFWNT9L_8tZ[348], b11_OFWNT9L_8tZ[347], 
        b11_OFWNT9L_8tZ[346], b11_OFWNT9L_8tZ[345], 
        b11_OFWNT9L_8tZ[344], b11_OFWNT9L_8tZ[343], 
        b11_OFWNT9L_8tZ[342], b11_OFWNT9L_8tZ[341], 
        b11_OFWNT9L_8tZ[340], b11_OFWNT9L_8tZ[339], 
        b11_OFWNT9L_8tZ[338], b11_OFWNT9L_8tZ[337], 
        b11_OFWNT9L_8tZ[336], b11_OFWNT9L_8tZ[335], 
        b11_OFWNT9L_8tZ[334], b11_OFWNT9L_8tZ[333], 
        b11_OFWNT9L_8tZ[332], b11_OFWNT9L_8tZ[331], 
        b11_OFWNT9L_8tZ[330], b11_OFWNT9L_8tZ[329], 
        b11_OFWNT9L_8tZ[328], b11_OFWNT9L_8tZ[327], 
        b11_OFWNT9L_8tZ[326], b11_OFWNT9L_8tZ[325], 
        b11_OFWNT9L_8tZ[324], b11_OFWNT9L_8tZ[323], 
        b11_OFWNT9L_8tZ[322], b11_OFWNT9L_8tZ[321], 
        b11_OFWNT9L_8tZ[320], b11_OFWNT9L_8tZ[319], 
        b11_OFWNT9L_8tZ[318], b11_OFWNT9L_8tZ[317], 
        b11_OFWNT9L_8tZ[316], b11_OFWNT9L_8tZ[315], 
        b11_OFWNT9L_8tZ[314], b11_OFWNT9L_8tZ[313], 
        b11_OFWNT9L_8tZ[312], b11_OFWNT9L_8tZ[311], 
        b11_OFWNT9L_8tZ[310], b11_OFWNT9L_8tZ[309], 
        b11_OFWNT9L_8tZ[308], b11_OFWNT9L_8tZ[307], 
        b11_OFWNT9L_8tZ[306], b11_OFWNT9L_8tZ[305], 
        b11_OFWNT9L_8tZ[304], b11_OFWNT9L_8tZ[303], 
        b11_OFWNT9L_8tZ[302], b11_OFWNT9L_8tZ[301], 
        b11_OFWNT9L_8tZ[300], b11_OFWNT9L_8tZ[299], 
        b11_OFWNT9L_8tZ[298], b11_OFWNT9L_8tZ[297], 
        b11_OFWNT9L_8tZ[296], b11_OFWNT9L_8tZ[295], 
        b11_OFWNT9L_8tZ[294], b11_OFWNT9L_8tZ[293], 
        b11_OFWNT9L_8tZ[292], b11_OFWNT9L_8tZ[291], 
        b11_OFWNT9L_8tZ[290], b11_OFWNT9L_8tZ[289], 
        b11_OFWNT9L_8tZ[288], b11_OFWNT9L_8tZ[287], 
        b11_OFWNT9L_8tZ[286], b11_OFWNT9L_8tZ[285], 
        b11_OFWNT9L_8tZ[284], b11_OFWNT9L_8tZ[283], 
        b11_OFWNT9L_8tZ[282], b11_OFWNT9L_8tZ[281], 
        b11_OFWNT9L_8tZ[280], b11_OFWNT9L_8tZ[279], 
        b11_OFWNT9L_8tZ[278], b11_OFWNT9L_8tZ[277], 
        b11_OFWNT9L_8tZ[276], b11_OFWNT9L_8tZ[275], 
        b11_OFWNT9L_8tZ[274], b11_OFWNT9L_8tZ[273], 
        b11_OFWNT9L_8tZ[272], b11_OFWNT9L_8tZ[271], 
        b11_OFWNT9L_8tZ[270], b11_OFWNT9L_8tZ[269], 
        b11_OFWNT9L_8tZ[268], b11_OFWNT9L_8tZ[267], 
        b11_OFWNT9L_8tZ[266], b11_OFWNT9L_8tZ[265], 
        b11_OFWNT9L_8tZ[264], b11_OFWNT9L_8tZ[263], 
        b11_OFWNT9L_8tZ[262], b11_OFWNT9L_8tZ[261], 
        b11_OFWNT9L_8tZ[260], b11_OFWNT9L_8tZ[259], 
        b11_OFWNT9L_8tZ[258], b11_OFWNT9L_8tZ[257], 
        b11_OFWNT9L_8tZ[256], b11_OFWNT9L_8tZ[255], 
        b11_OFWNT9L_8tZ[254], b11_OFWNT9L_8tZ[253], 
        b11_OFWNT9L_8tZ[252], b11_OFWNT9L_8tZ[251], 
        b11_OFWNT9L_8tZ[250], b11_OFWNT9L_8tZ[249], 
        b11_OFWNT9L_8tZ[248], b11_OFWNT9L_8tZ[247], 
        b11_OFWNT9L_8tZ[246], b11_OFWNT9L_8tZ[245], 
        b11_OFWNT9L_8tZ[244], b11_OFWNT9L_8tZ[243], 
        b11_OFWNT9L_8tZ[242], b11_OFWNT9L_8tZ[241], 
        b11_OFWNT9L_8tZ[240], b11_OFWNT9L_8tZ[239], 
        b11_OFWNT9L_8tZ[238], b11_OFWNT9L_8tZ[237], 
        b11_OFWNT9L_8tZ[236], b11_OFWNT9L_8tZ[235], 
        b11_OFWNT9L_8tZ[234], b11_OFWNT9L_8tZ[233], 
        b11_OFWNT9L_8tZ[232], b11_OFWNT9L_8tZ[231], 
        b11_OFWNT9L_8tZ[230], b11_OFWNT9L_8tZ[229], 
        b11_OFWNT9L_8tZ[228], b11_OFWNT9L_8tZ[227], 
        b11_OFWNT9L_8tZ[226], b11_OFWNT9L_8tZ[225], 
        b11_OFWNT9L_8tZ[224], b11_OFWNT9L_8tZ[223], 
        b11_OFWNT9L_8tZ[222], b11_OFWNT9L_8tZ[221], 
        b11_OFWNT9L_8tZ[220], b11_OFWNT9L_8tZ[219], 
        b11_OFWNT9L_8tZ[218], b11_OFWNT9L_8tZ[217], 
        b11_OFWNT9L_8tZ[216], b11_OFWNT9L_8tZ[215], 
        b11_OFWNT9L_8tZ[214], b11_OFWNT9L_8tZ[213], 
        b11_OFWNT9L_8tZ[212], b11_OFWNT9L_8tZ[211], 
        b11_OFWNT9L_8tZ[210], b11_OFWNT9L_8tZ[209], 
        b11_OFWNT9L_8tZ[208], b11_OFWNT9L_8tZ[207], 
        b11_OFWNT9L_8tZ[206], b11_OFWNT9L_8tZ[205], 
        b11_OFWNT9L_8tZ[204], b11_OFWNT9L_8tZ[203], 
        b11_OFWNT9L_8tZ[202], b11_OFWNT9L_8tZ[201], 
        b11_OFWNT9L_8tZ[200], b11_OFWNT9L_8tZ[199], 
        b11_OFWNT9L_8tZ[198], b11_OFWNT9L_8tZ[197], 
        b11_OFWNT9L_8tZ[196], b11_OFWNT9L_8tZ[195], 
        b11_OFWNT9L_8tZ[194], b11_OFWNT9L_8tZ[193], 
        b11_OFWNT9L_8tZ[192], b11_OFWNT9L_8tZ[191], 
        b11_OFWNT9L_8tZ[190], b11_OFWNT9L_8tZ[189], 
        b11_OFWNT9L_8tZ[188], b11_OFWNT9L_8tZ[187], 
        b11_OFWNT9L_8tZ[186], b11_OFWNT9L_8tZ[185], 
        b11_OFWNT9L_8tZ[184], b11_OFWNT9L_8tZ[183], 
        b11_OFWNT9L_8tZ[182], b11_OFWNT9L_8tZ[181], 
        b11_OFWNT9L_8tZ[180], b11_OFWNT9L_8tZ[179], 
        b11_OFWNT9L_8tZ[178], b11_OFWNT9L_8tZ[177], 
        b11_OFWNT9L_8tZ[176], b11_OFWNT9L_8tZ[175], 
        b11_OFWNT9L_8tZ[174], b11_OFWNT9L_8tZ[173], 
        b11_OFWNT9L_8tZ[172], b11_OFWNT9L_8tZ[171], 
        b11_OFWNT9L_8tZ[170], b11_OFWNT9L_8tZ[169], 
        b11_OFWNT9L_8tZ[168], b11_OFWNT9L_8tZ[167], 
        b11_OFWNT9L_8tZ[166], b11_OFWNT9L_8tZ[165], 
        b11_OFWNT9L_8tZ[164], b11_OFWNT9L_8tZ[163], 
        b11_OFWNT9L_8tZ[162], b11_OFWNT9L_8tZ[161], 
        b11_OFWNT9L_8tZ[160], b11_OFWNT9L_8tZ[159], 
        b11_OFWNT9L_8tZ[158], b11_OFWNT9L_8tZ[157], 
        b11_OFWNT9L_8tZ[156], b11_OFWNT9L_8tZ[155], 
        b11_OFWNT9L_8tZ[154], b11_OFWNT9L_8tZ[153], 
        b11_OFWNT9L_8tZ[152], b11_OFWNT9L_8tZ[151], 
        b11_OFWNT9L_8tZ[150], b11_OFWNT9L_8tZ[149], 
        b11_OFWNT9L_8tZ[148], b11_OFWNT9L_8tZ[147], 
        b11_OFWNT9L_8tZ[146], b11_OFWNT9L_8tZ[145], 
        b11_OFWNT9L_8tZ[144], b11_OFWNT9L_8tZ[143], 
        b11_OFWNT9L_8tZ[142], b11_OFWNT9L_8tZ[141], 
        b11_OFWNT9L_8tZ[140], b11_OFWNT9L_8tZ[139], 
        b11_OFWNT9L_8tZ[138], b11_OFWNT9L_8tZ[137], 
        b11_OFWNT9L_8tZ[136], b11_OFWNT9L_8tZ[135], 
        b11_OFWNT9L_8tZ[134], b11_OFWNT9L_8tZ[133], 
        b11_OFWNT9L_8tZ[132], b11_OFWNT9L_8tZ[131], 
        b11_OFWNT9L_8tZ[130], b11_OFWNT9L_8tZ[129], 
        b11_OFWNT9L_8tZ[128], b11_OFWNT9L_8tZ[127], 
        b11_OFWNT9L_8tZ[126], b11_OFWNT9L_8tZ[125], 
        b11_OFWNT9L_8tZ[124], b11_OFWNT9L_8tZ[123], 
        b11_OFWNT9L_8tZ[122], b11_OFWNT9L_8tZ[121], 
        b11_OFWNT9L_8tZ[120], b11_OFWNT9L_8tZ[119], 
        b11_OFWNT9L_8tZ[118], b11_OFWNT9L_8tZ[117], 
        b11_OFWNT9L_8tZ[116], b11_OFWNT9L_8tZ[115], 
        b11_OFWNT9L_8tZ[114], b11_OFWNT9L_8tZ[113], 
        b11_OFWNT9L_8tZ[112], b11_OFWNT9L_8tZ[111], 
        b11_OFWNT9L_8tZ[110], b11_OFWNT9L_8tZ[109], 
        b11_OFWNT9L_8tZ[108], b11_OFWNT9L_8tZ[107], 
        b11_OFWNT9L_8tZ[106], b11_OFWNT9L_8tZ[105], 
        b11_OFWNT9L_8tZ[104], b11_OFWNT9L_8tZ[103], 
        b11_OFWNT9L_8tZ[102], b11_OFWNT9L_8tZ[101], 
        b11_OFWNT9L_8tZ[100], b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], 
        b11_OFWNT9L_8tZ[97], b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], 
        b11_OFWNT9L_8tZ[94], b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], 
        b11_OFWNT9L_8tZ[91], b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], 
        b11_OFWNT9L_8tZ[88], b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], 
        b11_OFWNT9L_8tZ[85], b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], 
        b11_OFWNT9L_8tZ[82], b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], 
        b11_OFWNT9L_8tZ[79], b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], 
        b11_OFWNT9L_8tZ[76], b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], 
        b11_OFWNT9L_8tZ[73], b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], 
        b11_OFWNT9L_8tZ[70], b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], 
        b11_OFWNT9L_8tZ[67], b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], 
        b11_OFWNT9L_8tZ[64], b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], 
        b11_OFWNT9L_8tZ[61], b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], 
        b11_OFWNT9L_8tZ[58], b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], 
        b11_OFWNT9L_8tZ[55], b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], 
        b11_OFWNT9L_8tZ[52], b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], 
        b11_OFWNT9L_8tZ[49], b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], 
        b11_OFWNT9L_8tZ[46], b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], 
        b11_OFWNT9L_8tZ[43], b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], 
        b11_OFWNT9L_8tZ[40], b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], 
        b11_OFWNT9L_8tZ[37], b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], 
        b11_OFWNT9L_8tZ[34], b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], 
        b11_OFWNT9L_8tZ[31], b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], 
        b11_OFWNT9L_8tZ[28], b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], 
        b11_OFWNT9L_8tZ[25], b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], 
        b11_OFWNT9L_8tZ[22], b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], 
        b11_OFWNT9L_8tZ[19], b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], 
        b11_OFWNT9L_8tZ[16], b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], 
        b11_OFWNT9L_8tZ[13], b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], 
        b11_OFWNT9L_8tZ[10], b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], 
        b11_OFWNT9L_8tZ[7], b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], 
        b11_OFWNT9L_8tZ[4], b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], 
        b11_OFWNT9L_8tZ[1], b11_OFWNT9L_8tZ[0]}), .mdiclink_reg({
        mdiclink_reg[376], mdiclink_reg[375], mdiclink_reg[374], 
        mdiclink_reg[373], mdiclink_reg[372], mdiclink_reg[371], 
        mdiclink_reg[370], mdiclink_reg[369], mdiclink_reg[368], 
        mdiclink_reg[367], mdiclink_reg[366], mdiclink_reg[365], 
        mdiclink_reg[364], mdiclink_reg[363], mdiclink_reg[362], 
        mdiclink_reg[361], mdiclink_reg[360], mdiclink_reg[359], 
        mdiclink_reg[358], mdiclink_reg[357], mdiclink_reg[356], 
        mdiclink_reg[355], mdiclink_reg[354], mdiclink_reg[353], 
        mdiclink_reg[352], mdiclink_reg[351], mdiclink_reg[350], 
        mdiclink_reg[349], mdiclink_reg[348], mdiclink_reg[347], 
        mdiclink_reg[346], mdiclink_reg[345], mdiclink_reg[344], 
        mdiclink_reg[343], mdiclink_reg[342], mdiclink_reg[341], 
        mdiclink_reg[340], mdiclink_reg[339], mdiclink_reg[338], 
        mdiclink_reg[337], mdiclink_reg[336], mdiclink_reg[335], 
        mdiclink_reg[334], mdiclink_reg[333], mdiclink_reg[332], 
        mdiclink_reg[331], mdiclink_reg[330], mdiclink_reg[329], 
        mdiclink_reg[328], mdiclink_reg[327], mdiclink_reg[326], 
        mdiclink_reg[325], mdiclink_reg[324], mdiclink_reg[323], 
        mdiclink_reg[322], mdiclink_reg[321], mdiclink_reg[320], 
        mdiclink_reg[319], mdiclink_reg[318], mdiclink_reg[317], 
        mdiclink_reg[316], mdiclink_reg[315], mdiclink_reg[314], 
        mdiclink_reg[313], mdiclink_reg[312], mdiclink_reg[311], 
        mdiclink_reg[310], mdiclink_reg[309], mdiclink_reg[308], 
        mdiclink_reg[307], mdiclink_reg[306], mdiclink_reg[305], 
        mdiclink_reg[304], mdiclink_reg[303], mdiclink_reg[302], 
        mdiclink_reg[301], mdiclink_reg[300], mdiclink_reg[299], 
        mdiclink_reg[298], mdiclink_reg[297], mdiclink_reg[296], 
        mdiclink_reg[295], mdiclink_reg[294], mdiclink_reg[293], 
        mdiclink_reg[292], mdiclink_reg[291], mdiclink_reg[290], 
        mdiclink_reg[289], mdiclink_reg[288], mdiclink_reg[287], 
        mdiclink_reg[286], mdiclink_reg[285], mdiclink_reg[284], 
        mdiclink_reg[283], mdiclink_reg[282], mdiclink_reg[281], 
        mdiclink_reg[280], mdiclink_reg[279], mdiclink_reg[278], 
        mdiclink_reg[277], mdiclink_reg[276], mdiclink_reg[275], 
        mdiclink_reg[274], mdiclink_reg[273], mdiclink_reg[272], 
        mdiclink_reg[271], mdiclink_reg[270], mdiclink_reg[269], 
        mdiclink_reg[268], mdiclink_reg[267], mdiclink_reg[266], 
        mdiclink_reg[265], mdiclink_reg[264], mdiclink_reg[263], 
        mdiclink_reg[262], mdiclink_reg[261], mdiclink_reg[260], 
        mdiclink_reg[259], mdiclink_reg[258], mdiclink_reg[257], 
        mdiclink_reg[256], mdiclink_reg[255], mdiclink_reg[254], 
        mdiclink_reg[253], mdiclink_reg[252], mdiclink_reg[251], 
        mdiclink_reg[250], mdiclink_reg[249], mdiclink_reg[248], 
        mdiclink_reg[247], mdiclink_reg[246], mdiclink_reg[245], 
        mdiclink_reg[244], mdiclink_reg[243], mdiclink_reg[242], 
        mdiclink_reg[241], mdiclink_reg[240], mdiclink_reg[239], 
        mdiclink_reg[238], mdiclink_reg[237], mdiclink_reg[236], 
        mdiclink_reg[235], mdiclink_reg[234], mdiclink_reg[233], 
        mdiclink_reg[232], mdiclink_reg[231], mdiclink_reg[230], 
        mdiclink_reg[229], mdiclink_reg[228], mdiclink_reg[227], 
        mdiclink_reg[226], mdiclink_reg[225], mdiclink_reg[224], 
        mdiclink_reg[223], mdiclink_reg[222], mdiclink_reg[221], 
        mdiclink_reg[220], mdiclink_reg[219], mdiclink_reg[218], 
        mdiclink_reg[217], mdiclink_reg[216], mdiclink_reg[215], 
        mdiclink_reg[214], mdiclink_reg[213], mdiclink_reg[212], 
        mdiclink_reg[211], mdiclink_reg[210], mdiclink_reg[209], 
        mdiclink_reg[208], mdiclink_reg[207], mdiclink_reg[206], 
        mdiclink_reg[205], mdiclink_reg[204], mdiclink_reg[203], 
        mdiclink_reg[202], mdiclink_reg[201], mdiclink_reg[200], 
        mdiclink_reg[199], mdiclink_reg[198], mdiclink_reg[197], 
        mdiclink_reg[196], mdiclink_reg[195], mdiclink_reg[194], 
        mdiclink_reg[193], mdiclink_reg[192], mdiclink_reg[191], 
        mdiclink_reg[190], mdiclink_reg[189], mdiclink_reg[188], 
        mdiclink_reg[187], mdiclink_reg[186], mdiclink_reg[185], 
        mdiclink_reg[184], mdiclink_reg[183], mdiclink_reg[182], 
        mdiclink_reg[181], mdiclink_reg[180], mdiclink_reg[179], 
        mdiclink_reg[178], mdiclink_reg[177], mdiclink_reg[176], 
        mdiclink_reg[175], mdiclink_reg[174], mdiclink_reg[173], 
        mdiclink_reg[172], mdiclink_reg[171], mdiclink_reg[170], 
        mdiclink_reg[169], mdiclink_reg[168], mdiclink_reg[167], 
        mdiclink_reg[166], mdiclink_reg[165], mdiclink_reg[164], 
        mdiclink_reg[163], mdiclink_reg[162], mdiclink_reg[161], 
        mdiclink_reg[160], mdiclink_reg[159], mdiclink_reg[158], 
        mdiclink_reg[157], mdiclink_reg[156], mdiclink_reg[155], 
        mdiclink_reg[154], mdiclink_reg[153], mdiclink_reg[152], 
        mdiclink_reg[151], mdiclink_reg[150], mdiclink_reg[149], 
        mdiclink_reg[148], mdiclink_reg[147], mdiclink_reg[146], 
        mdiclink_reg[145], mdiclink_reg[144], mdiclink_reg[143], 
        mdiclink_reg[142], mdiclink_reg[141], mdiclink_reg[140], 
        mdiclink_reg[139], mdiclink_reg[138], mdiclink_reg[137], 
        mdiclink_reg[136], mdiclink_reg[135], mdiclink_reg[134], 
        mdiclink_reg[133], mdiclink_reg[132], mdiclink_reg[131], 
        mdiclink_reg[130], mdiclink_reg[129], mdiclink_reg[128], 
        mdiclink_reg[127], mdiclink_reg[126], mdiclink_reg[125], 
        mdiclink_reg[124], mdiclink_reg[123], mdiclink_reg[122], 
        mdiclink_reg[121], mdiclink_reg[120], mdiclink_reg[119], 
        mdiclink_reg[118], mdiclink_reg[117], mdiclink_reg[116], 
        mdiclink_reg[115], mdiclink_reg[114], mdiclink_reg[113], 
        mdiclink_reg[112], mdiclink_reg[111], mdiclink_reg[110], 
        mdiclink_reg[109], mdiclink_reg[108], mdiclink_reg[107], 
        mdiclink_reg[106], mdiclink_reg[105], mdiclink_reg[104], 
        mdiclink_reg[103], mdiclink_reg[102], mdiclink_reg[101], 
        mdiclink_reg[100], mdiclink_reg[99], mdiclink_reg[98], 
        mdiclink_reg[97], mdiclink_reg[96], mdiclink_reg[95], 
        mdiclink_reg[94], mdiclink_reg[93], mdiclink_reg[92], 
        mdiclink_reg[91], mdiclink_reg[90], mdiclink_reg[89], 
        mdiclink_reg[88], mdiclink_reg[87], mdiclink_reg[86], 
        mdiclink_reg[85], mdiclink_reg[84], mdiclink_reg[83], 
        mdiclink_reg[82], mdiclink_reg[81], mdiclink_reg[80], 
        mdiclink_reg[79], mdiclink_reg[78], mdiclink_reg[77], 
        mdiclink_reg[76], mdiclink_reg[75], mdiclink_reg[74], 
        mdiclink_reg[73], mdiclink_reg[72], mdiclink_reg[71], 
        mdiclink_reg[70], mdiclink_reg[69], mdiclink_reg[68], 
        mdiclink_reg[67], mdiclink_reg[66], mdiclink_reg[65], 
        mdiclink_reg[64], mdiclink_reg[63], mdiclink_reg[62], 
        mdiclink_reg[61], mdiclink_reg[60], mdiclink_reg[59], 
        mdiclink_reg[58], mdiclink_reg[57], mdiclink_reg[56], 
        mdiclink_reg[55], mdiclink_reg[54], mdiclink_reg[53], 
        mdiclink_reg[52], mdiclink_reg[51], mdiclink_reg[50], 
        mdiclink_reg[49], mdiclink_reg[48], mdiclink_reg[47], 
        mdiclink_reg[46], mdiclink_reg[45], mdiclink_reg[44], 
        mdiclink_reg[43], mdiclink_reg[42], mdiclink_reg[41], 
        mdiclink_reg[40], mdiclink_reg[39], mdiclink_reg[38], 
        mdiclink_reg[37], mdiclink_reg[36], mdiclink_reg[35], 
        mdiclink_reg[34], mdiclink_reg[33], mdiclink_reg[32], 
        mdiclink_reg[31], mdiclink_reg[30], mdiclink_reg[29], 
        mdiclink_reg[28], mdiclink_reg[27], mdiclink_reg[26], 
        mdiclink_reg[25], mdiclink_reg[24], mdiclink_reg[23], 
        mdiclink_reg[22], mdiclink_reg[21], mdiclink_reg[20], 
        mdiclink_reg[19], mdiclink_reg[18], mdiclink_reg[17], 
        mdiclink_reg[16], mdiclink_reg[15], mdiclink_reg[14], 
        mdiclink_reg[13], mdiclink_reg[12], mdiclink_reg[11], 
        mdiclink_reg[10], mdiclink_reg[9], mdiclink_reg[8], 
        mdiclink_reg[7], mdiclink_reg[6], mdiclink_reg[5], 
        mdiclink_reg[4], mdiclink_reg[3], mdiclink_reg[2], 
        mdiclink_reg[1], mdiclink_reg[0]}), .b6_Ocm0rW_0_0_o2({
        b6_Ocm0rW_0_0_o2[2]}), .b13_nAzGfFM_sLsv3({
        b13_nAzGfFM_sLsv3[1]}), .BW_clk_c(BW_clk_c), .b4_2o_z(b4_2o_z), 
        .b8_SoWGfWYY(b8_SoWGfWYY), .b13_oRB_MqCD2_EdR_RNI9OIA(
        b13_oRB_MqCD2_EdR_RNI9OIA));
    SLE \genblk9.b7_nYJ_BFM[168]  (.D(\b7_nYJ_BFM[167] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[168] ));
    SLE \genblk9.b7_nYJ_BFM[351]  (.D(\b7_nYJ_BFM[350] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[351] ));
    SLE \genblk9.b7_nYJ_BFM[148]  (.D(\b7_nYJ_BFM[147] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[148] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_168 (.A(\b7_nYJ_BFM[353] ), .B(
        \b7_nYJ_BFM[226] ), .C(\b7_vFW_PlM[352] ), .D(
        \b7_vFW_PlM[225] ), .Y(b3_PLF_168_net_1));
    SLE \genblk9.b7_nYJ_BFM[275]  (.D(\b7_nYJ_BFM[274] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[275] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_14 (.A(\b7_nYJ_BFM[147] ), .B(
        \b7_nYJ_BFM[20] ), .C(\b7_vFW_PlM[146] ), .D(\b7_vFW_PlM[19] ), 
        .Y(b3_PLF_14_net_1));
    SLE \genblk9.b7_nYJ_BFM[257]  (.D(\b7_nYJ_BFM[256] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[257] ));
    SLE \genblk9.b7_nYJ_BFM[76]  (.D(\b7_nYJ_BFM[75] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[76] ));
    SLE \genblk9.b7_nYJ_BFM[121]  (.D(\b7_nYJ_BFM[120] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[121] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_54 (.A(\b7_nYJ_BFM[286] ), .B(
        \b7_nYJ_BFM[30] ), .C(\b7_vFW_PlM[285] ), .D(\b7_vFW_PlM[29] ), 
        .Y(b3_PLF_54_net_1));
    SLE \genblk9.b7_nYJ_BFM[204]  (.D(\b7_nYJ_BFM[203] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[204] ));
    SLE \b12_PSyi_KyDbLbb[5]  (.D(\b12_2_St6KCa_jHv[5]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[5]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[137]  (.D(\b7_nYJ_BFM[136] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[137] ));
    SLE \genblk9.b7_nYJ_BFM[319]  (.D(\b7_nYJ_BFM[318] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[319] ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_76 (.A(\b7_nYJ_BFM[352] ), .B(
        \b7_nYJ_BFM[225] ), .C(\b7_vFW_PlM[351] ), .D(
        \b7_vFW_PlM[224] ), .Y(b3_PLF_76_net_1));
    SLE \genblk9.b7_nYJ_BFM[66]  (.D(\b7_nYJ_BFM[65] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[66] ));
    SLE \genblk9.b7_nYJ_BFM[41]  (.D(\b7_nYJ_BFM[40] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[41] ));
    SLE \genblk9.b7_nYJ_BFM[171]  (.D(\b7_nYJ_BFM[170] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[171] ));
    SLE \genblk9.b7_nYJ_BFM[215]  (.D(\b7_nYJ_BFM[214] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[215] ));
    SLE \genblk9.b7_nYJ_BFM[208]  (.D(\b7_nYJ_BFM[207] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[208] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_284 (.A(b3_PLF_8_net_1), .B(
        b3_PLF_7_net_1), .C(b3_PLF_6_net_1), .D(b3_PLF_5_net_1), .Y(
        b3_PLF_284_net_1));
    SLE \genblk9.b7_nYJ_BFM[82]  (.D(\b7_nYJ_BFM[81] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[82] ));
    SLE \b12_PSyi_KyDbLbb[8]  (.D(\b12_2_St6KCa_jHv[8]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[8]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[337]  (.D(\b7_nYJ_BFM[336] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[337] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_358 (.A(b3_PLF_304_net_1), .B(
        b3_PLF_303_net_1), .C(b3_PLF_302_net_1), .D(b3_PLF_301_net_1), 
        .Y(b3_PLF_358_net_1));
    SLE \genblk9.b7_nYJ_BFM[150]  (.D(\b7_nYJ_BFM[149] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[150] ));
    SLE \genblk9.b7_nYJ_BFM[338]  (.D(\b7_nYJ_BFM[337] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[338] ));
    SLE \genblk9.b7_nYJ_BFM[17]  (.D(\b7_nYJ_BFM[16] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[17] ));
    SLE \genblk9.b7_nYJ_BFM[109]  (.D(\b7_nYJ_BFM[108] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[109] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_311 (.A(b3_PLF_116_net_1), .B(
        b3_PLF_115_net_1), .C(b3_PLF_114_net_1), .D(b3_PLF_113_net_1), 
        .Y(b3_PLF_311_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_45 (.A(\b7_nYJ_BFM[330] ), .B(
        \b7_nYJ_BFM[74] ), .C(\b7_vFW_PlM[329] ), .D(\b7_vFW_PlM[73] ), 
        .Y(b3_PLF_45_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_295 (.A(b3_PLF_52_net_1), .B(
        b3_PLF_51_net_1), .C(b3_PLF_50_net_1), .D(b3_PLF_49_net_1), .Y(
        b3_PLF_295_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_315 (.A(b3_PLF_132_net_1), .B(
        b3_PLF_131_net_1), .C(b3_PLF_130_net_1), .D(b3_PLF_129_net_1), 
        .Y(b3_PLF_315_net_1));
    SLE \genblk9.b7_nYJ_BFM[299]  (.D(\b7_nYJ_BFM[298] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[299] ));
    SLE \genblk9.b7_nYJ_BFM[111]  (.D(\b7_nYJ_BFM[110] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[111] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_354 (.A(b3_PLF_288_net_1), .B(
        b3_PLF_287_net_1), .C(b3_PLF_286_net_1), .D(b3_PLF_285_net_1), 
        .Y(b3_PLF_354_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_48 (.A(\b7_nYJ_BFM[326] ), .B(
        \b7_nYJ_BFM[70] ), .C(\b7_vFW_PlM[325] ), .D(\b7_vFW_PlM[69] ), 
        .Y(b3_PLF_48_net_1));
    SLE \genblk9.b7_nYJ_BFM[23]  (.D(\b7_nYJ_BFM[22] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[23] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_127 (.A(\b7_nYJ_BFM[186] ), .B(
        \b7_nYJ_BFM[75] ), .C(\b7_vFW_PlM[185] ), .D(\b7_vFW_PlM[74] ), 
        .Y(b3_PLF_127_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_116 (.A(\b7_nYJ_BFM[297] ), .B(
        \b7_nYJ_BFM[170] ), .C(\b7_vFW_PlM[296] ), .D(
        \b7_vFW_PlM[169] ), .Y(b3_PLF_116_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[9]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_r_RNO_S[9] ), .Y(b9_v_mzCDYXs_3));
    SLE \genblk9.b7_nYJ_BFM[126]  (.D(\b7_nYJ_BFM[125] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[126] ));
    SLE \genblk9.b7_nYJ_BFM[96]  (.D(\b7_nYJ_BFM[95] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[96] ));
    CFG4 #( .INIT(16'hFEEE) )  b3_PLF_190 (.A(\un1_b4_BVmQ[1] ), .B(
        b3_PLF_4_net_1), .C(\b7_nYJ_BFM[258] ), .D(\b7_vFW_PlM[257] ), 
        .Y(b3_PLF_190_net_1));
    SLE \genblk9.b7_nYJ_BFM[300]  (.D(\b7_nYJ_BFM[299] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[300] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_2 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[2]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_1_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_2_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_2_net_1));
    SLE \genblk9.b7_nYJ_BFM[285]  (.D(\b7_nYJ_BFM[284] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[285] ));
    SLE \genblk9.b9_v_mzCDYXs[6]  (.D(b9_v_mzCDYXs_6), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[6] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_360 (.A(b3_PLF_312_net_1), .B(
        b3_PLF_311_net_1), .C(b3_PLF_310_net_1), .D(b3_PLF_309_net_1), 
        .Y(b3_PLF_360_net_1));
    SLE \genblk9.b7_nYJ_BFM[176]  (.D(\b7_nYJ_BFM[175] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[176] ));
    SLE \genblk9.b7_nYJ_BFM[262]  (.D(\b7_nYJ_BFM[261] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[262] ));
    SLE \genblk9.b7_nYJ_BFM[242]  (.D(\b7_nYJ_BFM[241] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[242] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_32 (.A(\b7_nYJ_BFM[331] ), .B(
        \b7_nYJ_BFM[203] ), .C(\b7_vFW_PlM[330] ), .D(
        \b7_vFW_PlM[202] ), .Y(b3_PLF_32_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_122 (.A(\b7_nYJ_BFM[289] ), .B(
        \b7_nYJ_BFM[162] ), .C(\b7_vFW_PlM[288] ), .D(
        \b7_vFW_PlM[161] ), .Y(b3_PLF_122_net_1));
    SLE \genblk9.b7_nYJ_BFM[105]  (.D(\b7_nYJ_BFM[104] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[105] ));
    SLE \genblk9.b7_nYJ_BFM[339]  (.D(\b7_nYJ_BFM[338] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[339] ));
    SLE \genblk9.b7_nYJ_BFM[103]  (.D(\b7_nYJ_BFM[102] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[103] ));
    SLE \genblk9.b7_nYJ_BFM[8]  (.D(\b7_nYJ_BFM[7] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[8] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_371 (.A(b3_PLF_356_net_1), .B(
        b3_PLF_355_net_1), .C(b3_PLF_354_net_1), .D(b3_PLF_353_net_1), 
        .Y(b3_PLF_371_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_158 (.A(\b7_nYJ_BFM[319] ), .B(
        \b7_nYJ_BFM[208] ), .C(\b7_vFW_PlM[318] ), .D(
        \b7_vFW_PlM[207] ), .Y(b3_PLF_158_net_1));
    SLE \genblk9.b7_nYJ_BFM[181]  (.D(\b7_nYJ_BFM[180] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[181] ));
    SLE \genblk9.b7_nYJ_BFM[235]  (.D(\b7_nYJ_BFM[234] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[235] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_363 (.A(b3_PLF_324_net_1), .B(
        b3_PLF_323_net_1), .C(b3_PLF_322_net_1), .D(b3_PLF_321_net_1), 
        .Y(b3_PLF_363_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_115 (.A(\b7_nYJ_BFM[76] ), .B(
        \b7_nYJ_BFM[59] ), .C(\b7_vFW_PlM[75] ), .D(\b7_vFW_PlM[58] ), 
        .Y(b3_PLF_115_net_1));
    SLE \genblk9.b7_nYJ_BFM[24]  (.D(\b7_nYJ_BFM[23] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[24] ));
    CFG3 #( .INIT(8'hF8) )  b3_PLF_188 (.A(\b7_nYJ_BFM[135] ), .B(
        \b7_vFW_PlM[134] ), .C(b3_PLF_0_net_1), .Y(b3_PLF_188_net_1));
    SLE \genblk9.b7_nYJ_BFM[116]  (.D(\b7_nYJ_BFM[115] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[116] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_176 (.A(\b7_nYJ_BFM[246] ), .B(
        \b7_nYJ_BFM[119] ), .C(\b7_vFW_PlM[245] ), .D(
        \b7_vFW_PlM[118] ), .Y(b3_PLF_176_net_1));
    SLE \genblk9.b7_nYJ_BFM[104]  (.D(\b7_nYJ_BFM[103] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[104] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_75 (.A(\b7_nYJ_BFM[354] ), .B(
        \b7_nYJ_BFM[98] ), .C(\b7_vFW_PlM[353] ), .D(\b7_vFW_PlM[97] ), 
        .Y(b3_PLF_75_net_1));
    SLE \genblk9.b7_nYJ_BFM[254]  (.D(\b7_nYJ_BFM[253] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[254] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_104 (.A(\b7_nYJ_BFM[154] ), .B(
        \b7_nYJ_BFM[43] ), .C(\b7_vFW_PlM[153] ), .D(\b7_vFW_PlM[42] ), 
        .Y(b3_PLF_104_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[5]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_5_S), .Y(b12_2_St6KCa_jHv_4));
    SLE \b12_2_St6KCa_jHv[7]  (.D(b12_2_St6KCa_jHv_6), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[7]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[131]  (.D(\b7_nYJ_BFM[130] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[131] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_78 (.A(\b7_nYJ_BFM[318] ), .B(
        \b7_nYJ_BFM[62] ), .C(\b7_vFW_PlM[317] ), .D(\b7_vFW_PlM[61] ), 
        .Y(b3_PLF_78_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_s_0_532 (.A(
        VCC_net_1), .B(b4_2o_z), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(un1_b12_2_St6KCa_jHv_s_0_532_FCO));
    SLE \b8_FZFFLXYE[1]  (.D(\b12_2_St6KCa_jHv[1]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[1]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[89]  (.D(\b7_nYJ_BFM[88] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[89] ));
    SLE \genblk9.b7_nYJ_BFM[77]  (.D(\b7_nYJ_BFM[76] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[77] ));
    SLE \genblk9.b7_nYJ_BFM[258]  (.D(\b7_nYJ_BFM[257] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[258] ));
    SLE \genblk9.b7_nYJ_BFM[50]  (.D(\b7_nYJ_BFM[49] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[50] ));
    SLE \genblk9.b7_nYJ_BFM[261]  (.D(\b7_nYJ_BFM[260] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[261] ));
    SLE \genblk9.b7_nYJ_BFM[241]  (.D(\b7_nYJ_BFM[240] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[241] ));
    SLE \genblk9.b7_nYJ_BFM[290]  (.D(\b7_nYJ_BFM[289] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[290] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_146 (.A(\b7_nYJ_BFM[192] ), .B(
        \b7_nYJ_BFM[65] ), .C(\b7_vFW_PlM[191] ), .D(\b7_vFW_PlM[64] ), 
        .Y(b3_PLF_146_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_175 (.A(\b7_nYJ_BFM[375] ), .B(
        \b7_nYJ_BFM[248] ), .C(\b7_vFW_PlM[374] ), .D(
        \b7_vFW_PlM[247] ), .Y(b3_PLF_175_net_1));
    SLE \genblk9.b7_nYJ_BFM[30]  (.D(\b7_nYJ_BFM[29] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[30] ));
    SLE \genblk9.b7_nYJ_BFM[186]  (.D(\b7_nYJ_BFM[185] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[186] ));
    SLE \genblk9.b7_nYJ_BFM[67]  (.D(\b7_nYJ_BFM[66] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[67] ));
    SLE \genblk9.b7_nYJ_BFM[159]  (.D(\b7_nYJ_BFM[158] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[159] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_134 (.A(\b7_nYJ_BFM[305] ), .B(
        \b7_nYJ_BFM[49] ), .C(\b7_vFW_PlM[304] ), .D(\b7_vFW_PlM[48] ), 
        .Y(b3_PLF_134_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_80 (.A(\b7_nYJ_BFM[267] ), .B(
        \b7_nYJ_BFM[28] ), .C(\b7_vFW_PlM[266] ), .D(\b7_vFW_PlM[27] ), 
        .Y(b3_PLF_80_net_1));
    CFG4 #( .INIT(16'h2000) )  b7_yYh03wy_u_0_a2 (.A(IICE_comm2iice_0), 
        .B(IICE_comm2iice_4), .C(b7_yYh03wy_u_0_m2_net_1), .D(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .Y(b7_yYh03wy));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_111 (.A(\b7_nYJ_BFM[273] ), .B(
        \b7_nYJ_BFM[17] ), .C(\b7_vFW_PlM[272] ), .D(\b7_vFW_PlM[16] ), 
        .Y(b3_PLF_111_net_1));
    SLE \genblk9.b7_nYJ_BFM[203]  (.D(\b7_nYJ_BFM[202] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[203] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_60 (.A(\b7_nYJ_BFM[342] ), .B(
        \b7_nYJ_BFM[86] ), .C(\b7_vFW_PlM[341] ), .D(\b7_vFW_PlM[85] ), 
        .Y(b3_PLF_60_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_289 (.A(b3_PLF_28_net_1), .B(
        b3_PLF_27_net_1), .C(b3_PLF_26_net_1), .D(b3_PLF_25_net_1), .Y(
        b3_PLF_289_net_1));
    SLE \genblk9.b7_nYJ_BFM[102]  (.D(\b7_nYJ_BFM[101] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[102] ));
    SLE \genblk9.b7_nYJ_BFM[350]  (.D(\b7_nYJ_BFM[349] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[350] ));
    SLE \b8_FZFFLXYE[9]  (.D(\b12_2_St6KCa_jHv[9]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[9]_net_1 ));
    SLE \b8_FZFFLXYE[5]  (.D(\b12_2_St6KCa_jHv[5]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[5]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_19 (.A(\b7_nYJ_BFM[204] ), .B(
        \b7_nYJ_BFM[93] ), .C(\b7_vFW_PlM[203] ), .D(\b7_vFW_PlM[92] ), 
        .Y(b3_PLF_19_net_1));
    SLE \genblk9.b7_nYJ_BFM[136]  (.D(\b7_nYJ_BFM[135] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[136] ));
    SLE \genblk9.b7_nYJ_BFM[325]  (.D(\b7_nYJ_BFM[324] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[325] ));
    SLE \genblk9.b7_nYJ_BFM[88]  (.D(\b7_nYJ_BFM[87] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[88] ));
    SLE \genblk9.b7_nYJ_BFM[363]  (.D(\b7_nYJ_BFM[362] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[363] ));
    SLE \genblk9.b7_nYJ_BFM[343]  (.D(\b7_nYJ_BFM[342] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[343] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_145 (.A(\b7_nYJ_BFM[321] ), .B(
        \b7_nYJ_BFM[194] ), .C(\b7_vFW_PlM[320] ), .D(
        \b7_vFW_PlM[193] ), .Y(b3_PLF_145_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_83 (.A(\b7_nYJ_BFM[247] ), .B(
        \b7_nYJ_BFM[120] ), .C(\b7_vFW_PlM[246] ), .D(
        \b7_vFW_PlM[119] ), .Y(b3_PLF_83_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_59 (.A(\b7_nYJ_BFM[215] ), .B(
        \b7_nYJ_BFM[88] ), .C(\b7_vFW_PlM[214] ), .D(\b7_vFW_PlM[87] ), 
        .Y(b3_PLF_59_net_1));
    SLE \genblk9.b7_nYJ_BFM[229]  (.D(\b7_nYJ_BFM[228] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[229] ));
    SLE \genblk9.b7_nYJ_BFM[155]  (.D(\b7_nYJ_BFM[154] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[155] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_63 (.A(\b7_nYJ_BFM[338] ), .B(
        \b7_nYJ_BFM[82] ), .C(\b7_vFW_PlM[337] ), .D(\b7_vFW_PlM[81] ), 
        .Y(b3_PLF_63_net_1));
    SLE \genblk9.b7_nYJ_BFM[97]  (.D(\b7_nYJ_BFM[96] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[97] ));
    SLE \genblk9.b7_nYJ_BFM[42]  (.D(\b7_nYJ_BFM[41] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[42] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_160 (.A(\b7_nYJ_BFM[285] ), .B(
        \b7_nYJ_BFM[29] ), .C(\b7_vFW_PlM[284] ), .D(\b7_vFW_PlM[28] ), 
        .Y(b3_PLF_160_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_353 (.A(b3_PLF_187_net_1), .B(
        b3_PLF_281_net_1), .C(b3_PLF_188_net_1), .D(b3_PLF_330_net_1), 
        .Y(b3_PLF_353_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_163 (.A(\b7_nYJ_BFM[232] ), .B(
        \b7_nYJ_BFM[105] ), .C(\b7_vFW_PlM[231] ), .D(
        \b7_vFW_PlM[104] ), .Y(b3_PLF_163_net_1));
    SLE \genblk9.b7_nYJ_BFM[153]  (.D(\b7_nYJ_BFM[152] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[153] ));
    SLE \genblk9.b7_nYJ_BFM[375]  (.D(\b7_nYJ_BFM[374] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[375] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_171 (.A(\b7_nYJ_BFM[301] ), .B(
        \b7_nYJ_BFM[190] ), .C(\b7_vFW_PlM[300] ), .D(
        \b7_vFW_PlM[189] ), .Y(b3_PLF_171_net_1));
    SLE \genblk9.b7_nYJ_BFM[279]  (.D(\b7_nYJ_BFM[278] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[279] ));
    SLE \genblk9.b7_nYJ_BFM[15]  (.D(\b7_nYJ_BFM[14] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[15] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_119 (.A(\b7_nYJ_BFM[293] ), .B(
        \b7_nYJ_BFM[166] ), .C(\b7_vFW_PlM[292] ), .D(
        \b7_vFW_PlM[165] ), .Y(b3_PLF_119_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_292 (.A(b3_PLF_40_net_1), .B(
        b3_PLF_39_net_1), .C(b3_PLF_38_net_1), .D(b3_PLF_37_net_1), .Y(
        b3_PLF_292_net_1));
    SLE \genblk9.b7_nYJ_BFM[266]  (.D(\b7_nYJ_BFM[265] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[266] ));
    SLE \genblk9.b7_nYJ_BFM[246]  (.D(\b7_nYJ_BFM[245] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[246] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIQD3J7[8]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[8] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_7), .S(\b9_v_mzCDYXs_RNIQD3J7_S[8] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_8));
    SLE \genblk9.b7_nYJ_BFM[154]  (.D(\b7_nYJ_BFM[153] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[154] ));
    SLE \genblk9.b7_nYJ_BFM[26]  (.D(\b7_nYJ_BFM[25] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[26] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_319 (.A(b3_PLF_148_net_1), .B(
        b3_PLF_147_net_1), .C(b3_PLF_146_net_1), .D(b3_PLF_145_net_1), 
        .Y(b3_PLF_319_net_1));
    SLE \genblk9.b7_nYJ_BFM[315]  (.D(\b7_nYJ_BFM[314] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[315] ));
    SLE \genblk9.b7_nYJ_BFM[219]  (.D(\b7_nYJ_BFM[218] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[219] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_91 (.A(\b7_nYJ_BFM[300] ), .B(
        \b7_nYJ_BFM[189] ), .C(\b7_vFW_PlM[299] ), .D(
        \b7_vFW_PlM[188] ), .Y(b3_PLF_91_net_1));
    SLE \genblk9.b7_nYJ_BFM[297]  (.D(\b7_nYJ_BFM[296] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[297] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_316 (.A(b3_PLF_136_net_1), .B(
        b3_PLF_135_net_1), .C(b3_PLF_134_net_1), .D(b3_PLF_133_net_1), 
        .Y(b3_PLF_316_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_5 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[5]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_4_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_5_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_5_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_141 (.A(\b7_nYJ_BFM[327] ), .B(
        \b7_nYJ_BFM[71] ), .C(\b7_vFW_PlM[326] ), .D(\b7_vFW_PlM[70] ), 
        .Y(b3_PLF_141_net_1));
    SLE \genblk9.b7_nYJ_BFM[108]  (.D(\b7_nYJ_BFM[107] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[108] ));
    CFG2 #( .INIT(4'h8) )  \genblk9.un1_b4_BVmQ[1]  (.A(
        \b7_vFW_PlM[1] ), .B(\b7_nYJ_BFM[2] ), .Y(\un1_b4_BVmQ[1] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[1]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNIA2R45_S[1] ), .Y(b9_v_mzCDYXs_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_179 (.A(\b7_nYJ_BFM[242] ), .B(
        \b7_nYJ_BFM[115] ), .C(\b7_vFW_PlM[241] ), .D(
        \b7_vFW_PlM[114] ), .Y(b3_PLF_179_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_124 (.A(\b7_nYJ_BFM[366] ), .B(
        \b7_nYJ_BFM[271] ), .C(\b7_vFW_PlM[365] ), .D(
        \b7_vFW_PlM[270] ), .Y(b3_PLF_124_net_1));
    SLE \genblk9.b7_nYJ_BFM[326]  (.D(\b7_nYJ_BFM[325] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[326] ));
    SLE \genblk9.b7_nYJ_BFM[253]  (.D(\b7_nYJ_BFM[252] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[253] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_308 (.A(b3_PLF_104_net_1), .B(
        b3_PLF_103_net_1), .C(b3_PLF_102_net_1), .D(b3_PLF_101_net_1), 
        .Y(b3_PLF_308_net_1));
    SLE \genblk9.b7_nYJ_BFM[53]  (.D(\b7_nYJ_BFM[52] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[53] ));
    SLE \genblk9.b7_nYJ_BFM[11]  (.D(\b7_nYJ_BFM[10] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[11] ));
    CFG4 #( .INIT(16'h8000) )  b8_jAA_KlCO_0_sqmuxa_8 (.A(
        \b12_2_St6KCa_jHv[7]_net_1 ), .B(b8_jAA_KlCO_0_sqmuxa_6_net_1), 
        .C(b4_2o_z), .D(\b12_2_St6KCa_jHv[8]_net_1 ), .Y(
        b8_jAA_KlCO_0_sqmuxa_8_net_1));
    SLE \genblk9.b7_nYJ_BFM[9]  (.D(\b7_nYJ_BFM[8] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[9] ));
    SLE \genblk9.b7_nYJ_BFM[190]  (.D(\b7_nYJ_BFM[189] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[190] ));
    SLE \b12_2_St6KCa_jHv[2]  (.D(b12_2_St6KCa_jHv_1), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[2]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[152]  (.D(\b7_nYJ_BFM[151] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[152] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_40 (.A(\b7_nYJ_BFM[304] ), .B(
        \b7_nYJ_BFM[177] ), .C(\b7_vFW_PlM[303] ), .D(
        \b7_vFW_PlM[176] ), .Y(b3_PLF_40_net_1));
    SLE \genblk9.b7_nYJ_BFM[220]  (.D(\b7_nYJ_BFM[219] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[220] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_297 (.A(b3_PLF_60_net_1), .B(
        b3_PLF_59_net_1), .C(b3_PLF_58_net_1), .D(b3_PLF_57_net_1), .Y(
        b3_PLF_297_net_1));
    SLE \genblk9.b7_nYJ_BFM[289]  (.D(\b7_nYJ_BFM[288] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[289] ));
    SLE \genblk9.b7_nYJ_BFM[33]  (.D(\b7_nYJ_BFM[32] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[33] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_357 (.A(b3_PLF_300_net_1), .B(
        b3_PLF_299_net_1), .C(b3_PLF_298_net_1), .D(b3_PLF_297_net_1), 
        .Y(b3_PLF_357_net_1));
    SLE \genblk9.b7_nYJ_BFM[376]  (.D(\b7_nYJ_BFM[375] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[376] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_304 (.A(b3_PLF_88_net_1), .B(
        b3_PLF_87_net_1), .C(b3_PLF_86_net_1), .D(b3_PLF_85_net_1), .Y(
        b3_PLF_304_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_285 (.A(b3_PLF_12_net_1), .B(
        b3_PLF_11_net_1), .C(b3_PLF_10_net_1), .D(b3_PLF_9_net_1), .Y(
        b3_PLF_285_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_97 (.A(\b7_nYJ_BFM[132] ), .B(
        \b7_nYJ_BFM[5] ), .C(\b7_vFW_PlM[131] ), .D(\b7_vFW_PlM[4] ), 
        .Y(b3_PLF_97_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[2]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI95U74[383] ), .C(
        \b9_v_mzCDYXs_RNINN0G5_S[2] ), .Y(b9_v_mzCDYXs_0));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_150 (.A(\b7_nYJ_BFM[218] ), .B(
        \b7_nYJ_BFM[107] ), .C(\b7_vFW_PlM[217] ), .D(
        \b7_vFW_PlM[106] ), .Y(b3_PLF_150_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[2]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_2_S), .Y(b12_2_St6KCa_jHv_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_153 (.A(\b7_nYJ_BFM[214] ), .B(
        \b7_nYJ_BFM[87] ), .C(\b7_vFW_PlM[213] ), .D(\b7_vFW_PlM[86] ), 
        .Y(b3_PLF_153_net_1));
    SLE \genblk9.b7_nYJ_BFM[270]  (.D(\b7_nYJ_BFM[269] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[270] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_82 (.A(\b7_nYJ_BFM[376] ), .B(
        \b7_nYJ_BFM[249] ), .C(\b7_vFW_PlM[375] ), .D(
        \b7_vFW_PlM[248] ), .Y(b3_PLF_82_net_1));
    SLE \genblk9.b7_nYJ_BFM[49]  (.D(\b7_nYJ_BFM[48] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[49] ));
    SLE \genblk9.b7_nYJ_BFM[324]  (.D(\b7_nYJ_BFM[323] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[324] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_180 (.A(\b7_nYJ_BFM[369] ), .B(
        \b7_nYJ_BFM[113] ), .C(\b7_vFW_PlM[368] ), .D(
        \b7_vFW_PlM[112] ), .Y(b3_PLF_180_net_1));
    SLE \genblk9.b7_nYJ_BFM[75]  (.D(\b7_nYJ_BFM[74] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[75] ));
    SLE \genblk9.b7_nYJ_BFM[335]  (.D(\b7_nYJ_BFM[334] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[335] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_62 (.A(\b7_nYJ_BFM[211] ), .B(
        \b7_nYJ_BFM[84] ), .C(\b7_vFW_PlM[210] ), .D(\b7_vFW_PlM[83] ), 
        .Y(b3_PLF_62_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_293 (.A(b3_PLF_44_net_1), .B(
        b3_PLF_43_net_1), .C(b3_PLF_42_net_1), .D(b3_PLF_41_net_1), .Y(
        b3_PLF_293_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_149 (.A(\b7_nYJ_BFM[364] ), .B(
        \b7_nYJ_BFM[124] ), .C(\b7_vFW_PlM[363] ), .D(
        \b7_vFW_PlM[123] ), .Y(b3_PLF_149_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_302 (.A(b3_PLF_80_net_1), .B(
        b3_PLF_79_net_1), .C(b3_PLF_78_net_1), .D(b3_PLF_77_net_1), .Y(
        b3_PLF_302_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_21 (.A(\b7_nYJ_BFM[298] ), .B(
        \b7_nYJ_BFM[42] ), .C(\b7_vFW_PlM[297] ), .D(\b7_vFW_PlM[41] ), 
        .Y(b3_PLF_21_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_183 (.A(\b7_nYJ_BFM[317] ), .B(
        \b7_nYJ_BFM[61] ), .C(\b7_vFW_PlM[316] ), .D(\b7_vFW_PlM[60] ), 
        .Y(b3_PLF_183_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_16 (.A(\b7_nYJ_BFM[272] ), .B(
        \b7_nYJ_BFM[145] ), .C(\b7_vFW_PlM[271] ), .D(
        \b7_vFW_PlM[144] ), .Y(b3_PLF_16_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_8 (.A(\b7_nYJ_BFM[299] ), .B(
        \b7_nYJ_BFM[171] ), .C(\b7_vFW_PlM[298] ), .D(
        \b7_vFW_PlM[170] ), .Y(b3_PLF_8_net_1));
    SLE \genblk9.b7_nYJ_BFM[239]  (.D(\b7_nYJ_BFM[238] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[239] ));
    SLE \genblk9.b7_nYJ_BFM[316]  (.D(\b7_nYJ_BFM[315] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[316] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_6 (.A(\b7_nYJ_BFM[333] ), .B(
        \b7_nYJ_BFM[222] ), .C(\b7_vFW_PlM[332] ), .D(
        \b7_vFW_PlM[221] ), .Y(b3_PLF_6_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_43 (.A(\b7_nYJ_BFM[236] ), .B(
        \b7_nYJ_BFM[125] ), .C(\b7_vFW_PlM[235] ), .D(
        \b7_vFW_PlM[124] ), .Y(b3_PLF_43_net_1));
    SLE \genblk9.b7_nYJ_BFM[54]  (.D(\b7_nYJ_BFM[53] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[54] ));
    SLE \genblk9.b7_nYJ_BFM[65]  (.D(\b7_nYJ_BFM[64] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[65] ));
    SLE \genblk9.b7_nYJ_BFM[374]  (.D(\b7_nYJ_BFM[373] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[7] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[374] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_56 (.A(\b7_nYJ_BFM[363] ), .B(
        \b7_nYJ_BFM[235] ), .C(\b7_vFW_PlM[362] ), .D(
        \b7_vFW_PlM[234] ), .Y(b3_PLF_56_net_1));
    SLE \b12_2_St6KCa_jHv[1]  (.D(b12_2_St6KCa_jHv_0), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[1]_net_1 ));
    
endmodule


module b7_PLF_6lN_x_0(
       b13_nvmFL_fx2rbuQ,
       b16_nYhI39swMeEd_A78,
       b12_vABZ3qsY_Lyh,
       b7_yYh03wy,
       b13_nUTQBgfDb_Z4D,
       N_8,
       b3_PLF_sn_N_12,
       b11_vABZ3qsY_XH_2,
       b3_PLF_sn_N_17,
       b15_OFWNT9khWqH_R9k,
       b12_uRrc2XfY_Lyh,
       b3_PLF_u_d_bm,
       b13_PSyiBgfDb_Z4D,
       b3_PLF_u_d_am
    );
input  [6:1] b13_nvmFL_fx2rbuQ;
input  b16_nYhI39swMeEd_A78;
input  b12_vABZ3qsY_Lyh;
input  b7_yYh03wy;
input  b13_nUTQBgfDb_Z4D;
output N_8;
output b3_PLF_sn_N_12;
output b11_vABZ3qsY_XH_2;
output b3_PLF_sn_N_17;
input  b15_OFWNT9khWqH_R9k;
input  b12_uRrc2XfY_Lyh;
output b3_PLF_u_d_bm;
input  b13_PSyiBgfDb_Z4D;
output b3_PLF_u_d_am;

    wire b3_PLF_sn_N_20, N_6, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hC0A0) )  b3_PLF_u_d_bm_inst_1 (.A(
        b15_OFWNT9khWqH_R9k), .B(b12_uRrc2XfY_Lyh), .C(
        b11_vABZ3qsY_XH_2), .D(b13_nvmFL_fx2rbuQ[3]), .Y(b3_PLF_u_d_bm)
        );
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hD8) )  b3_PLF_4 (.A(b13_nvmFL_fx2rbuQ[6]), .B(
        b7_yYh03wy), .C(b13_nUTQBgfDb_Z4D), .Y(N_8));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h88D8) )  b3_PLF_u_d_am_inst_1 (.A(
        b13_nvmFL_fx2rbuQ[3]), .B(N_6), .C(b13_PSyiBgfDb_Z4D), .D(
        b13_nvmFL_fx2rbuQ[2]), .Y(b3_PLF_u_d_am));
    CFG3 #( .INIT(8'h01) )  b3_PLF_6_0 (.A(b13_nvmFL_fx2rbuQ[4]), .B(
        b13_nvmFL_fx2rbuQ[6]), .C(b13_nvmFL_fx2rbuQ[5]), .Y(
        b11_vABZ3qsY_XH_2));
    CFG4 #( .INIT(16'h5FFE) )  b3_PLF_sn_m16 (.A(b13_nvmFL_fx2rbuQ[6]), 
        .B(b3_PLF_sn_N_20), .C(b13_nvmFL_fx2rbuQ[5]), .D(
        b13_nvmFL_fx2rbuQ[4]), .Y(b3_PLF_sn_N_17));
    CFG2 #( .INIT(4'h4) )  b3_PLF_sn_m14_e (.A(b13_nvmFL_fx2rbuQ[1]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .Y(b3_PLF_sn_N_20));
    CFG3 #( .INIT(8'h4E) )  b3_PLF_sn_m11 (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[1]), .C(b13_nvmFL_fx2rbuQ[2]), .Y(
        b3_PLF_sn_N_12));
    CFG3 #( .INIT(8'hE4) )  b3_PLF_0 (.A(b13_nvmFL_fx2rbuQ[1]), .B(
        b16_nYhI39swMeEd_A78), .C(b12_vABZ3qsY_Lyh), .Y(N_6));
    
endmodule


module b12_nvmFL_la1xyH_x_0(
       b13_nvmFL_fx2rbuQ,
       b11_vABZ3qsY_XH_2,
       b11_uRrc_9urXBb,
       b12_PSyiBgfDb_bd,
       b3_PLF_sn_N_17,
       b3_PLF_u_d_bm,
       b3_PLF,
       b3_PLF_sn_N_12,
       b3_PLF_u_d_am,
       N_8,
       b14_OFWNT9khWqH_3i,
       b15_nYhI39swMeEd_Mg,
       b12_nUTQBgfDb_bd,
       b11_vABZ3qsY_XH,
       b12_ibScJX_E2_bd,
       b12_PSyi2XfYF_bd,
       b11_uRrc2XfY_XH
    );
input  [6:1] b13_nvmFL_fx2rbuQ;
input  b11_vABZ3qsY_XH_2;
input  b11_uRrc_9urXBb;
output b12_PSyiBgfDb_bd;
input  b3_PLF_sn_N_17;
input  b3_PLF_u_d_bm;
output b3_PLF;
input  b3_PLF_sn_N_12;
input  b3_PLF_u_d_am;
input  N_8;
output b14_OFWNT9khWqH_3i;
output b15_nYhI39swMeEd_Mg;
output b12_nUTQBgfDb_bd;
output b11_vABZ3qsY_XH;
output b12_ibScJX_E2_bd;
output b12_PSyi2XfYF_bd;
output b11_uRrc2XfY_XH;

    wire b9_nvmFLR_ab_2, b3_PLF_1_net_1, b9_nvmFLz_ab_1, 
        b9_nvmFLp_ab_1, b9_nvmFLm_ab_2_net_1, b9_nvmFLm_ab_3_net_1, 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h2000) )  b9_nvmFLT_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .C(b9_nvmFLp_ab_1), .D(
        b11_vABZ3qsY_XH_2), .Y(b11_vABZ3qsY_XH));
    CFG4 #( .INIT(16'h1000) )  b9_nvmFLH_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[1]), .C(b11_vABZ3qsY_XH_2), .D(
        b9_nvmFLz_ab_1), .Y(b14_OFWNT9khWqH_3i));
    CFG2 #( .INIT(4'h1) )  b9_nvmFLm_ab_2 (.A(b13_nvmFL_fx2rbuQ[1]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .Y(b9_nvmFLm_ab_2_net_1));
    CFG4 #( .INIT(16'h4000) )  b9_nvmFLp_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .C(b11_vABZ3qsY_XH_2), .D(
        b9_nvmFLp_ab_1), .Y(b12_PSyi2XfYF_bd));
    CFG4 #( .INIT(16'h04BF) )  b3_PLF_1 (.A(b13_nvmFL_fx2rbuQ[6]), .B(
        b3_PLF_sn_N_12), .C(b3_PLF_u_d_am), .D(N_8), .Y(b3_PLF_1_net_1)
        );
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hA202) )  b3_PLF_inst_1 (.A(b11_uRrc_9urXBb), .B(
        b3_PLF_1_net_1), .C(b3_PLF_sn_N_17), .D(b3_PLF_u_d_bm), .Y(
        b3_PLF));
    CFG2 #( .INIT(4'h8) )  b9_nvmFLR_ab_1 (.A(b11_uRrc_9urXBb), .B(
        b13_nvmFL_fx2rbuQ[1]), .Y(b9_nvmFLp_ab_1));
    CFG4 #( .INIT(16'h2000) )  b9_nvmFLm_ab_3 (.A(b13_nvmFL_fx2rbuQ[4])
        , .B(b13_nvmFL_fx2rbuQ[3]), .C(b11_uRrc_9urXBb), .D(
        b9_nvmFLm_ab_2_net_1), .Y(b9_nvmFLm_ab_3_net_1));
    CFG4 #( .INIT(16'h2000) )  b9_nvmFLz_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[1]), .C(b11_vABZ3qsY_XH_2), .D(
        b9_nvmFLz_ab_1), .Y(b11_uRrc2XfY_XH));
    CFG3 #( .INIT(8'h10) )  b9_nvmFLm_ab (.A(b13_nvmFL_fx2rbuQ[6]), .B(
        b13_nvmFL_fx2rbuQ[5]), .C(b9_nvmFLm_ab_3_net_1), .Y(
        b12_ibScJX_E2_bd));
    CFG4 #( .INIT(16'h8000) )  b9_nvmFLP_ab0 (.A(b11_vABZ3qsY_XH_2), 
        .B(b11_uRrc_9urXBb), .C(b13_nvmFL_fx2rbuQ[3]), .D(
        b9_nvmFLm_ab_2_net_1), .Y(b15_nYhI39swMeEd_Mg));
    CFG4 #( .INIT(16'h0800) )  b9_nvmFLQ_ab (.A(b11_vABZ3qsY_XH_2), .B(
        b11_uRrc_9urXBb), .C(b13_nvmFL_fx2rbuQ[1]), .D(b9_nvmFLR_ab_2), 
        .Y(b12_nUTQBgfDb_bd));
    CFG4 #( .INIT(16'h8000) )  b9_nvmFLR_ab (.A(b11_vABZ3qsY_XH_2), .B(
        b11_uRrc_9urXBb), .C(b13_nvmFL_fx2rbuQ[1]), .D(b9_nvmFLR_ab_2), 
        .Y(b12_PSyiBgfDb_bd));
    CFG2 #( .INIT(4'h1) )  b9_nvmFLQ_ab_2 (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .Y(b9_nvmFLR_ab_2));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  b9_nvmFLH_ab_1 (.A(b11_uRrc_9urXBb), .B(
        b13_nvmFL_fx2rbuQ[2]), .Y(b9_nvmFLz_ab_1));
    
endmodule


module b3_uKr_x(
       b13_nvmFL_fx2rbuQ,
       b11_uRrc_9urXBb,
       b3_PLy,
       b3_PLF,
       b7_PLy_PlM,
       b12_PSyiBgfDb_bd,
       b12_PSyi2XfYF_bd,
       b14_OFWNT9khWqH_3i,
       b13_PSyiBgfDb_Z4D,
       b13_PSyi2XfYF_Z4D,
       b15_OFWNT9khWqH_R9k,
       b7_yYh03wy,
       b12_nUTQBgfDb_bd,
       b11_uRrc2XfY_XH,
       b13_nUTQBgfDb_Z4D,
       b15_nYhI39swMeEd_Mg,
       b16_nYhI39swMeEd_A78,
       b11_vABZ3qsY_XH,
       b12_vABZ3qsY_Lyh,
       b12_ibScJX_E2_bd,
       b13_ibScJX_E2_Z4D,
       b12_uRrc2XfY_Lyh
    );
input  [6:1] b13_nvmFL_fx2rbuQ;
input  b11_uRrc_9urXBb;
input  b3_PLy;
output b3_PLF;
output b7_PLy_PlM;
output b12_PSyiBgfDb_bd;
output b12_PSyi2XfYF_bd;
output b14_OFWNT9khWqH_3i;
input  b13_PSyiBgfDb_Z4D;
input  b13_PSyi2XfYF_Z4D;
input  b15_OFWNT9khWqH_R9k;
input  b7_yYh03wy;
output b12_nUTQBgfDb_bd;
output b11_uRrc2XfY_XH;
input  b13_nUTQBgfDb_Z4D;
output b15_nYhI39swMeEd_Mg;
input  b16_nYhI39swMeEd_A78;
output b11_vABZ3qsY_XH;
input  b12_vABZ3qsY_Lyh;
output b12_ibScJX_E2_bd;
input  b13_ibScJX_E2_Z4D;
input  b12_uRrc2XfY_Lyh;

    wire b3_PLy_net_1, GND_net_1, VCC_net_1, 
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_12 , 
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_17 , N_8, b11_vABZ3qsY_XH_2, 
        b3_PLF_u_d_am, b3_PLF_u_d_bm;
    assign b3_PLy_net_1 = b3_PLy;
    assign b7_PLy_PlM = b3_PLy_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    b7_PLF_6lN_x_0 b12_PLF_6lN_8tYv (.b13_nvmFL_fx2rbuQ({
        b13_nvmFL_fx2rbuQ[6], b13_nvmFL_fx2rbuQ[5], 
        b13_nvmFL_fx2rbuQ[4], b13_nvmFL_fx2rbuQ[3], 
        b13_nvmFL_fx2rbuQ[2], b13_nvmFL_fx2rbuQ[1]}), 
        .b16_nYhI39swMeEd_A78(b16_nYhI39swMeEd_A78), .b12_vABZ3qsY_Lyh(
        b12_vABZ3qsY_Lyh), .b7_yYh03wy(b7_yYh03wy), .b13_nUTQBgfDb_Z4D(
        b13_nUTQBgfDb_Z4D), .N_8(N_8), .b3_PLF_sn_N_12(
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_12 ), .b11_vABZ3qsY_XH_2(
        b11_vABZ3qsY_XH_2), .b3_PLF_sn_N_17(
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_17 ), .b15_OFWNT9khWqH_R9k(
        b15_OFWNT9khWqH_R9k), .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh), 
        .b3_PLF_u_d_bm(b3_PLF_u_d_bm), .b13_PSyiBgfDb_Z4D(
        b13_PSyiBgfDb_Z4D), .b3_PLF_u_d_am(b3_PLF_u_d_am));
    b12_nvmFL_la1xyH_x_0 b10_nvscB_rGsL (.b13_nvmFL_fx2rbuQ({
        b13_nvmFL_fx2rbuQ[6], b13_nvmFL_fx2rbuQ[5], 
        b13_nvmFL_fx2rbuQ[4], b13_nvmFL_fx2rbuQ[3], 
        b13_nvmFL_fx2rbuQ[2], b13_nvmFL_fx2rbuQ[1]}), 
        .b11_vABZ3qsY_XH_2(b11_vABZ3qsY_XH_2), .b11_uRrc_9urXBb(
        b11_uRrc_9urXBb), .b12_PSyiBgfDb_bd(b12_PSyiBgfDb_bd), 
        .b3_PLF_sn_N_17(\b12_PLF_6lN_8tYv.b3_PLF_sn_N_17 ), 
        .b3_PLF_u_d_bm(b3_PLF_u_d_bm), .b3_PLF(b3_PLF), 
        .b3_PLF_sn_N_12(\b12_PLF_6lN_8tYv.b3_PLF_sn_N_12 ), 
        .b3_PLF_u_d_am(b3_PLF_u_d_am), .N_8(N_8), .b14_OFWNT9khWqH_3i(
        b14_OFWNT9khWqH_3i), .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), 
        .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), .b11_vABZ3qsY_XH(
        b11_vABZ3qsY_XH), .b12_ibScJX_E2_bd(b12_ibScJX_E2_bd), 
        .b12_PSyi2XfYF_bd(b12_PSyi2XfYF_bd), .b11_uRrc2XfY_XH(
        b11_uRrc2XfY_XH));
    
endmodule


module IICE_x(
       BW_c,
       BW_out_c,
       dac_count,
       dac1_db_c,
       \data_from_adc[8] ,
       \data_from_adc[7] ,
       \data_from_adc[6] ,
       \data_from_adc[4] ,
       \data_from_adc[5] ,
       \data_from_adc[3] ,
       \data_from_adc[2] ,
       \data_from_adc[1] ,
       \data_from_adc[0] ,
       fpga_count,
       fr_adc_count,
       fpga_shift_2,
       sdv_count,
       temp1,
       temp2,
       temp3,
       temp_count_data,
       temp_count,
       dds_sin,
       dds_cos,
       IICE_comm2iice,
       freq_2,
       freq_14,
       freq_15,
       freq_0,
       freq_1,
       freq_6,
       freq_10,
       freq_11,
       freq_13,
       BW_clk_c,
       clk_dac2,
       dac1_clk_c,
       temp_sck_c,
       temp1_csn_c,
       temp2_csn_c,
       temp3_csn_c,
       temp_so_c,
       IICE_iice2comm
    );
input  [14:0] BW_c;
input  [14:0] BW_out_c;
input  [7:1] dac_count;
input  [13:5] dac1_db_c;
input  [11:0] \data_from_adc[8] ;
input  [11:0] \data_from_adc[7] ;
input  [11:0] \data_from_adc[6] ;
input  [11:0] \data_from_adc[4] ;
input  [11:0] \data_from_adc[5] ;
input  [11:0] \data_from_adc[3] ;
input  [11:0] \data_from_adc[2] ;
input  [11:0] \data_from_adc[1] ;
input  [11:0] \data_from_adc[0] ;
input  [14:0] fpga_count;
input  [3:1] fr_adc_count;
input  [14:0] fpga_shift_2;
input  [1:0] sdv_count;
input  [15:0] temp1;
input  [15:0] temp2;
input  [15:0] temp3;
input  [4:0] temp_count_data;
input  [31:0] temp_count;
input  [7:0] dds_sin;
input  [7:0] dds_cos;
input  [11:0] IICE_comm2iice;
input  freq_2;
input  freq_14;
input  freq_15;
input  freq_0;
input  freq_1;
input  freq_6;
input  freq_10;
input  freq_11;
input  freq_13;
input  BW_clk_c;
input  clk_dac2;
input  dac1_clk_c;
input  temp_sck_c;
input  temp1_csn_c;
input  temp2_csn_c;
input  temp3_csn_c;
input  temp_so_c;
output IICE_iice2comm;

    wire \mdiclink_reg[6]_net_1 , VCC_net_1, GND_net_1, 
        \mdiclink_reg[5]_net_1 , \mdiclink_reg[4]_net_1 , 
        \mdiclink_reg[3]_net_1 , \mdiclink_reg[2]_net_1 , 
        \mdiclink_reg[1]_net_1 , \mdiclink_reg[0]_net_1 , 
        \mdiclink_reg[21]_net_1 , \mdiclink_reg[20]_net_1 , 
        \mdiclink_reg[19]_net_1 , \mdiclink_reg[18]_net_1 , 
        \mdiclink_reg[17]_net_1 , \mdiclink_reg[16]_net_1 , 
        \mdiclink_reg[15]_net_1 , \mdiclink_reg[14]_net_1 , 
        \mdiclink_reg[13]_net_1 , \mdiclink_reg[12]_net_1 , 
        \mdiclink_reg[11]_net_1 , \mdiclink_reg[10]_net_1 , 
        \mdiclink_reg[9]_net_1 , \mdiclink_reg[8]_net_1 , 
        \mdiclink_reg[7]_net_1 , \mdiclink_reg[36]_net_1 , 
        \mdiclink_reg[35]_net_1 , \mdiclink_reg[34]_net_1 , 
        \mdiclink_reg[33]_net_1 , \mdiclink_reg[32]_net_1 , 
        \mdiclink_reg[31]_net_1 , \mdiclink_reg[30]_net_1 , 
        \mdiclink_reg[29]_net_1 , \mdiclink_reg[28]_net_1 , 
        \mdiclink_reg[27]_net_1 , \mdiclink_reg[26]_net_1 , 
        \mdiclink_reg[25]_net_1 , \mdiclink_reg[24]_net_1 , 
        \mdiclink_reg[23]_net_1 , \mdiclink_reg[22]_net_1 , 
        \mdiclink_reg[51]_net_1 , \mdiclink_reg[50]_net_1 , 
        \mdiclink_reg[49]_net_1 , \mdiclink_reg[48]_net_1 , 
        \mdiclink_reg[47]_net_1 , \mdiclink_reg[46]_net_1 , 
        \mdiclink_reg[45]_net_1 , \mdiclink_reg[44]_net_1 , 
        \mdiclink_reg[43]_net_1 , \mdiclink_reg[42]_net_1 , 
        \mdiclink_reg[41]_net_1 , \mdiclink_reg[40]_net_1 , 
        \mdiclink_reg[39]_net_1 , \mdiclink_reg[38]_net_1 , 
        \mdiclink_reg[37]_net_1 , \mdiclink_reg[66]_net_1 , 
        \mdiclink_reg[65]_net_1 , \mdiclink_reg[64]_net_1 , 
        \mdiclink_reg[63]_net_1 , \mdiclink_reg[62]_net_1 , 
        \mdiclink_reg[61]_net_1 , \mdiclink_reg[60]_net_1 , 
        \mdiclink_reg[59]_net_1 , \mdiclink_reg[58]_net_1 , 
        \mdiclink_reg[57]_net_1 , \mdiclink_reg[56]_net_1 , 
        \mdiclink_reg[55]_net_1 , \mdiclink_reg[54]_net_1 , 
        \mdiclink_reg[53]_net_1 , \mdiclink_reg[52]_net_1 , 
        \mdiclink_reg[81]_net_1 , \mdiclink_reg[80]_net_1 , 
        \mdiclink_reg[79]_net_1 , \mdiclink_reg[78]_net_1 , 
        \mdiclink_reg[77]_net_1 , \mdiclink_reg[76]_net_1 , 
        \mdiclink_reg[75]_net_1 , \mdiclink_reg[74]_net_1 , 
        \mdiclink_reg[73]_net_1 , \mdiclink_reg[72]_net_1 , 
        \mdiclink_reg[71]_net_1 , \mdiclink_reg[70]_net_1 , 
        \mdiclink_reg[69]_net_1 , \mdiclink_reg[68]_net_1 , 
        \mdiclink_reg[67]_net_1 , \mdiclink_reg[96]_net_1 , 
        \mdiclink_reg[95]_net_1 , \mdiclink_reg[94]_net_1 , 
        \mdiclink_reg[93]_net_1 , \mdiclink_reg[92]_net_1 , 
        \mdiclink_reg[91]_net_1 , \mdiclink_reg[90]_net_1 , 
        \mdiclink_reg[89]_net_1 , \mdiclink_reg[88]_net_1 , 
        \mdiclink_reg[87]_net_1 , \mdiclink_reg[86]_net_1 , 
        \mdiclink_reg[85]_net_1 , \mdiclink_reg[84]_net_1 , 
        \mdiclink_reg[83]_net_1 , \mdiclink_reg[82]_net_1 , 
        \mdiclink_reg[111]_net_1 , \mdiclink_reg[110]_net_1 , 
        \mdiclink_reg[109]_net_1 , \mdiclink_reg[108]_net_1 , 
        \mdiclink_reg[107]_net_1 , \mdiclink_reg[106]_net_1 , 
        \mdiclink_reg[105]_net_1 , \mdiclink_reg[104]_net_1 , 
        \mdiclink_reg[103]_net_1 , \mdiclink_reg[102]_net_1 , 
        \mdiclink_reg[101]_net_1 , \mdiclink_reg[100]_net_1 , 
        \mdiclink_reg[99]_net_1 , \mdiclink_reg[98]_net_1 , 
        \mdiclink_reg[97]_net_1 , \mdiclink_reg[126]_net_1 , 
        \mdiclink_reg[125]_net_1 , \mdiclink_reg[124]_net_1 , 
        \mdiclink_reg[123]_net_1 , \mdiclink_reg[122]_net_1 , 
        \mdiclink_reg[121]_net_1 , \mdiclink_reg[120]_net_1 , 
        \mdiclink_reg[119]_net_1 , \mdiclink_reg[118]_net_1 , 
        \mdiclink_reg[117]_net_1 , \mdiclink_reg[116]_net_1 , 
        \mdiclink_reg[115]_net_1 , \mdiclink_reg[114]_net_1 , 
        \mdiclink_reg[113]_net_1 , \mdiclink_reg[112]_net_1 , 
        \mdiclink_reg[141]_net_1 , \mdiclink_reg[140]_net_1 , 
        \mdiclink_reg[139]_net_1 , \mdiclink_reg[138]_net_1 , 
        \mdiclink_reg[137]_net_1 , \mdiclink_reg[136]_net_1 , 
        \mdiclink_reg[135]_net_1 , \mdiclink_reg[134]_net_1 , 
        \mdiclink_reg[133]_net_1 , \mdiclink_reg[132]_net_1 , 
        \mdiclink_reg[131]_net_1 , \mdiclink_reg[130]_net_1 , 
        \mdiclink_reg[129]_net_1 , \mdiclink_reg[128]_net_1 , 
        \mdiclink_reg[127]_net_1 , \mdiclink_reg[156]_net_1 , 
        \mdiclink_reg[155]_net_1 , \mdiclink_reg[154]_net_1 , 
        \mdiclink_reg[153]_net_1 , \mdiclink_reg[152]_net_1 , 
        \mdiclink_reg[151]_net_1 , \mdiclink_reg[150]_net_1 , 
        \mdiclink_reg[149]_net_1 , \mdiclink_reg[148]_net_1 , 
        \mdiclink_reg[147]_net_1 , \mdiclink_reg[146]_net_1 , 
        \mdiclink_reg[145]_net_1 , \mdiclink_reg[144]_net_1 , 
        \mdiclink_reg[143]_net_1 , \mdiclink_reg[142]_net_1 , 
        \mdiclink_reg[157]_net_1 , \mdiclink_reg[186]_net_1 , 
        \mdiclink_reg[185]_net_1 , \mdiclink_reg[184]_net_1 , 
        \mdiclink_reg[183]_net_1 , \mdiclink_reg[182]_net_1 , 
        \mdiclink_reg[181]_net_1 , \mdiclink_reg[180]_net_1 , 
        \mdiclink_reg[179]_net_1 , \mdiclink_reg[178]_net_1 , 
        \mdiclink_reg[177]_net_1 , \mdiclink_reg[176]_net_1 , 
        \mdiclink_reg[175]_net_1 , \mdiclink_reg[174]_net_1 , 
        \mdiclink_reg[201]_net_1 , \mdiclink_reg[200]_net_1 , 
        \mdiclink_reg[199]_net_1 , \mdiclink_reg[198]_net_1 , 
        \mdiclink_reg[197]_net_1 , \mdiclink_reg[196]_net_1 , 
        \mdiclink_reg[195]_net_1 , \mdiclink_reg[194]_net_1 , 
        \mdiclink_reg[193]_net_1 , \mdiclink_reg[192]_net_1 , 
        \mdiclink_reg[191]_net_1 , \mdiclink_reg[190]_net_1 , 
        \mdiclink_reg[189]_net_1 , \mdiclink_reg[188]_net_1 , 
        \mdiclink_reg[187]_net_1 , \mdiclink_reg[216]_net_1 , 
        \mdiclink_reg[215]_net_1 , \mdiclink_reg[214]_net_1 , 
        \mdiclink_reg[213]_net_1 , \mdiclink_reg[212]_net_1 , 
        \mdiclink_reg[211]_net_1 , \mdiclink_reg[210]_net_1 , 
        \mdiclink_reg[209]_net_1 , \mdiclink_reg[208]_net_1 , 
        \mdiclink_reg[207]_net_1 , \mdiclink_reg[206]_net_1 , 
        \mdiclink_reg[205]_net_1 , \mdiclink_reg[204]_net_1 , 
        \mdiclink_reg[203]_net_1 , \mdiclink_reg[202]_net_1 , 
        \mdiclink_reg[231]_net_1 , \mdiclink_reg[230]_net_1 , 
        \mdiclink_reg[229]_net_1 , \mdiclink_reg[228]_net_1 , 
        \mdiclink_reg[227]_net_1 , \mdiclink_reg[226]_net_1 , 
        \mdiclink_reg[225]_net_1 , \mdiclink_reg[224]_net_1 , 
        \mdiclink_reg[223]_net_1 , \mdiclink_reg[222]_net_1 , 
        \mdiclink_reg[221]_net_1 , \mdiclink_reg[220]_net_1 , 
        \mdiclink_reg[219]_net_1 , \mdiclink_reg[218]_net_1 , 
        \mdiclink_reg[217]_net_1 , \mdiclink_reg[246]_net_1 , 
        \mdiclink_reg[245]_net_1 , \mdiclink_reg[244]_net_1 , 
        \mdiclink_reg[243]_net_1 , \mdiclink_reg[242]_net_1 , 
        \mdiclink_reg[241]_net_1 , \mdiclink_reg[240]_net_1 , 
        \mdiclink_reg[239]_net_1 , \mdiclink_reg[238]_net_1 , 
        \mdiclink_reg[237]_net_1 , \mdiclink_reg[236]_net_1 , 
        \mdiclink_reg[235]_net_1 , \mdiclink_reg[234]_net_1 , 
        \mdiclink_reg[233]_net_1 , \mdiclink_reg[232]_net_1 , 
        \mdiclink_reg[261]_net_1 , \mdiclink_reg[260]_net_1 , 
        \mdiclink_reg[259]_net_1 , \mdiclink_reg[258]_net_1 , 
        \mdiclink_reg[257]_net_1 , \mdiclink_reg[256]_net_1 , 
        \mdiclink_reg[255]_net_1 , \mdiclink_reg[254]_net_1 , 
        \mdiclink_reg[253]_net_1 , \mdiclink_reg[252]_net_1 , 
        \mdiclink_reg[251]_net_1 , \mdiclink_reg[250]_net_1 , 
        \mdiclink_reg[249]_net_1 , \mdiclink_reg[248]_net_1 , 
        \mdiclink_reg[247]_net_1 , \mdiclink_reg[276]_net_1 , 
        \mdiclink_reg[275]_net_1 , \mdiclink_reg[274]_net_1 , 
        \mdiclink_reg[273]_net_1 , \mdiclink_reg[272]_net_1 , 
        \mdiclink_reg[271]_net_1 , \mdiclink_reg[270]_net_1 , 
        \mdiclink_reg[269]_net_1 , \mdiclink_reg[268]_net_1 , 
        \mdiclink_reg[267]_net_1 , \mdiclink_reg[266]_net_1 , 
        \mdiclink_reg[265]_net_1 , \mdiclink_reg[264]_net_1 , 
        \mdiclink_reg[263]_net_1 , \mdiclink_reg[262]_net_1 , 
        \mdiclink_reg[291]_net_1 , \mdiclink_reg[290]_net_1 , 
        \mdiclink_reg[289]_net_1 , \mdiclink_reg[288]_net_1 , 
        \mdiclink_reg[287]_net_1 , \mdiclink_reg[286]_net_1 , 
        \mdiclink_reg[285]_net_1 , \mdiclink_reg[284]_net_1 , 
        \mdiclink_reg[283]_net_1 , \mdiclink_reg[282]_net_1 , 
        \mdiclink_reg[281]_net_1 , \mdiclink_reg[280]_net_1 , 
        \mdiclink_reg[279]_net_1 , \mdiclink_reg[278]_net_1 , 
        \mdiclink_reg[277]_net_1 , \mdiclink_reg[306]_net_1 , 
        \mdiclink_reg[305]_net_1 , \mdiclink_reg[304]_net_1 , 
        \mdiclink_reg[303]_net_1 , \mdiclink_reg[302]_net_1 , 
        \mdiclink_reg[301]_net_1 , \mdiclink_reg[300]_net_1 , 
        \mdiclink_reg[299]_net_1 , \mdiclink_reg[298]_net_1 , 
        \mdiclink_reg[297]_net_1 , \mdiclink_reg[296]_net_1 , 
        \mdiclink_reg[295]_net_1 , \mdiclink_reg[294]_net_1 , 
        \mdiclink_reg[293]_net_1 , \mdiclink_reg[292]_net_1 , 
        \mdiclink_reg[321]_net_1 , \mdiclink_reg[320]_net_1 , 
        \mdiclink_reg[319]_net_1 , \mdiclink_reg[318]_net_1 , 
        \mdiclink_reg[317]_net_1 , \mdiclink_reg[316]_net_1 , 
        \mdiclink_reg[315]_net_1 , \mdiclink_reg[314]_net_1 , 
        \mdiclink_reg[313]_net_1 , \mdiclink_reg[312]_net_1 , 
        \mdiclink_reg[311]_net_1 , \mdiclink_reg[310]_net_1 , 
        \mdiclink_reg[309]_net_1 , \mdiclink_reg[308]_net_1 , 
        \mdiclink_reg[307]_net_1 , \mdiclink_reg[336]_net_1 , 
        \mdiclink_reg[335]_net_1 , \mdiclink_reg[334]_net_1 , 
        \mdiclink_reg[333]_net_1 , \mdiclink_reg[332]_net_1 , 
        \mdiclink_reg[331]_net_1 , \mdiclink_reg[330]_net_1 , 
        \mdiclink_reg[329]_net_1 , \mdiclink_reg[328]_net_1 , 
        \mdiclink_reg[327]_net_1 , \mdiclink_reg[326]_net_1 , 
        \mdiclink_reg[325]_net_1 , \mdiclink_reg[324]_net_1 , 
        \mdiclink_reg[323]_net_1 , \mdiclink_reg[322]_net_1 , 
        \mdiclink_reg[351]_net_1 , \mdiclink_reg[350]_net_1 , 
        \mdiclink_reg[349]_net_1 , \mdiclink_reg[348]_net_1 , 
        \mdiclink_reg[347]_net_1 , \mdiclink_reg[346]_net_1 , 
        \mdiclink_reg[345]_net_1 , \mdiclink_reg[344]_net_1 , 
        \mdiclink_reg[343]_net_1 , \mdiclink_reg[342]_net_1 , 
        \mdiclink_reg[341]_net_1 , \mdiclink_reg[340]_net_1 , 
        \mdiclink_reg[339]_net_1 , \mdiclink_reg[338]_net_1 , 
        \mdiclink_reg[337]_net_1 , \mdiclink_reg[366]_net_1 , 
        \mdiclink_reg[365]_net_1 , \mdiclink_reg[364]_net_1 , 
        \mdiclink_reg[363]_net_1 , \mdiclink_reg[362]_net_1 , 
        \mdiclink_reg[361]_net_1 , \mdiclink_reg[360]_net_1 , 
        \mdiclink_reg[359]_net_1 , \mdiclink_reg[358]_net_1 , 
        \mdiclink_reg[357]_net_1 , \mdiclink_reg[356]_net_1 , 
        \mdiclink_reg[355]_net_1 , \mdiclink_reg[354]_net_1 , 
        \mdiclink_reg[353]_net_1 , \mdiclink_reg[352]_net_1 , 
        \mdiclink_reg[376]_net_1 , \mdiclink_reg[375]_net_1 , 
        \mdiclink_reg[374]_net_1 , \mdiclink_reg[373]_net_1 , 
        \mdiclink_reg[372]_net_1 , \mdiclink_reg[371]_net_1 , 
        \mdiclink_reg[370]_net_1 , \mdiclink_reg[369]_net_1 , 
        \mdiclink_reg[368]_net_1 , \mdiclink_reg[367]_net_1 , 
        \mdiclink_reg[158]_net_1 , \mdiclink_reg[173]_net_1 , 
        \mdiclink_reg[172]_net_1 , \mdiclink_reg[171]_net_1 , 
        \mdiclink_reg[170]_net_1 , \mdiclink_reg[169]_net_1 , 
        \mdiclink_reg[168]_net_1 , \mdiclink_reg[167]_net_1 , 
        \mdiclink_reg[166]_net_1 , \mdiclink_reg[165]_net_1 , 
        \mdiclink_reg[164]_net_1 , \mdiclink_reg[163]_net_1 , 
        \mdiclink_reg[162]_net_1 , \mdiclink_reg[161]_net_1 , 
        \mdiclink_reg[160]_net_1 , \mdiclink_reg[159]_net_1 , b4_PLyF, 
        b8_PSyiBgYG, b8_PSyi2XYG, b10_OFWNT9khFt, b7_PSyi3wy, 
        b9_OFWNT9Mxf, b7_yYh03wy, b12_nUTQBgfDb_bd, b11_uRrc2XfY_XH, 
        b13_nUTQBgfDb_Z4D, b15_nYhI39swMeEd_Mg, b16_nYhI39swMeEd_A78, 
        b11_vABZ3qsY_XH, b12_vABZ3qsY_Lyh, b12_ibScJX_E2_bd, 
        b12_uRrc2XfY_Lyh, \b6_Ocm0rW_0_0_o2[2] , 
        \b13_nAzGfFM_sLsv3[1] , \b11_OFWNT9L_8tZ[0] , 
        \b11_OFWNT9L_8tZ[1] , \b11_OFWNT9L_8tZ[2] , 
        \b11_OFWNT9L_8tZ[3] , \b11_OFWNT9L_8tZ[4] , 
        \b11_OFWNT9L_8tZ[5] , \b11_OFWNT9L_8tZ[6] , 
        \b11_OFWNT9L_8tZ[7] , \b11_OFWNT9L_8tZ[8] , 
        \b11_OFWNT9L_8tZ[9] , \b11_OFWNT9L_8tZ[10] , 
        \b11_OFWNT9L_8tZ[11] , \b11_OFWNT9L_8tZ[12] , 
        \b11_OFWNT9L_8tZ[13] , \b11_OFWNT9L_8tZ[14] , 
        \b11_OFWNT9L_8tZ[15] , \b11_OFWNT9L_8tZ[16] , 
        \b11_OFWNT9L_8tZ[17] , \b11_OFWNT9L_8tZ[18] , 
        \b11_OFWNT9L_8tZ[19] , \b11_OFWNT9L_8tZ[20] , 
        \b11_OFWNT9L_8tZ[21] , \b11_OFWNT9L_8tZ[22] , 
        \b11_OFWNT9L_8tZ[23] , \b11_OFWNT9L_8tZ[24] , 
        \b11_OFWNT9L_8tZ[25] , \b11_OFWNT9L_8tZ[26] , 
        \b11_OFWNT9L_8tZ[27] , \b11_OFWNT9L_8tZ[28] , 
        \b11_OFWNT9L_8tZ[29] , \b11_OFWNT9L_8tZ[30] , 
        \b11_OFWNT9L_8tZ[31] , \b11_OFWNT9L_8tZ[32] , 
        \b11_OFWNT9L_8tZ[33] , \b11_OFWNT9L_8tZ[34] , 
        \b11_OFWNT9L_8tZ[35] , \b11_OFWNT9L_8tZ[36] , 
        \b11_OFWNT9L_8tZ[37] , \b11_OFWNT9L_8tZ[38] , 
        \b11_OFWNT9L_8tZ[39] , \b11_OFWNT9L_8tZ[40] , 
        \b11_OFWNT9L_8tZ[41] , \b11_OFWNT9L_8tZ[42] , 
        \b11_OFWNT9L_8tZ[43] , \b11_OFWNT9L_8tZ[44] , 
        \b11_OFWNT9L_8tZ[45] , \b11_OFWNT9L_8tZ[46] , 
        \b11_OFWNT9L_8tZ[47] , \b11_OFWNT9L_8tZ[48] , 
        \b11_OFWNT9L_8tZ[49] , \b11_OFWNT9L_8tZ[50] , 
        \b11_OFWNT9L_8tZ[51] , \b11_OFWNT9L_8tZ[52] , 
        \b11_OFWNT9L_8tZ[53] , \b11_OFWNT9L_8tZ[54] , 
        \b11_OFWNT9L_8tZ[55] , \b11_OFWNT9L_8tZ[56] , 
        \b11_OFWNT9L_8tZ[57] , \b11_OFWNT9L_8tZ[58] , 
        \b11_OFWNT9L_8tZ[59] , \b11_OFWNT9L_8tZ[60] , 
        \b11_OFWNT9L_8tZ[61] , \b11_OFWNT9L_8tZ[62] , 
        \b11_OFWNT9L_8tZ[63] , \b11_OFWNT9L_8tZ[64] , 
        \b11_OFWNT9L_8tZ[65] , \b11_OFWNT9L_8tZ[66] , 
        \b11_OFWNT9L_8tZ[67] , \b11_OFWNT9L_8tZ[68] , 
        \b11_OFWNT9L_8tZ[69] , \b11_OFWNT9L_8tZ[70] , 
        \b11_OFWNT9L_8tZ[71] , \b11_OFWNT9L_8tZ[72] , 
        \b11_OFWNT9L_8tZ[73] , \b11_OFWNT9L_8tZ[74] , 
        \b11_OFWNT9L_8tZ[75] , \b11_OFWNT9L_8tZ[76] , 
        \b11_OFWNT9L_8tZ[77] , \b11_OFWNT9L_8tZ[78] , 
        \b11_OFWNT9L_8tZ[79] , \b11_OFWNT9L_8tZ[80] , 
        \b11_OFWNT9L_8tZ[81] , \b11_OFWNT9L_8tZ[82] , 
        \b11_OFWNT9L_8tZ[83] , \b11_OFWNT9L_8tZ[84] , 
        \b11_OFWNT9L_8tZ[85] , \b11_OFWNT9L_8tZ[86] , 
        \b11_OFWNT9L_8tZ[87] , \b11_OFWNT9L_8tZ[88] , 
        \b11_OFWNT9L_8tZ[89] , \b11_OFWNT9L_8tZ[90] , 
        \b11_OFWNT9L_8tZ[91] , \b11_OFWNT9L_8tZ[92] , 
        \b11_OFWNT9L_8tZ[93] , \b11_OFWNT9L_8tZ[94] , 
        \b11_OFWNT9L_8tZ[95] , \b11_OFWNT9L_8tZ[96] , 
        \b11_OFWNT9L_8tZ[97] , \b11_OFWNT9L_8tZ[98] , 
        \b11_OFWNT9L_8tZ[99] , \b11_OFWNT9L_8tZ[100] , 
        \b11_OFWNT9L_8tZ[101] , \b11_OFWNT9L_8tZ[102] , 
        \b11_OFWNT9L_8tZ[103] , \b11_OFWNT9L_8tZ[104] , 
        \b11_OFWNT9L_8tZ[105] , \b11_OFWNT9L_8tZ[106] , 
        \b11_OFWNT9L_8tZ[107] , \b11_OFWNT9L_8tZ[108] , 
        \b11_OFWNT9L_8tZ[109] , \b11_OFWNT9L_8tZ[110] , 
        \b11_OFWNT9L_8tZ[111] , \b11_OFWNT9L_8tZ[112] , 
        \b11_OFWNT9L_8tZ[113] , \b11_OFWNT9L_8tZ[114] , 
        \b11_OFWNT9L_8tZ[115] , \b11_OFWNT9L_8tZ[116] , 
        \b11_OFWNT9L_8tZ[117] , \b11_OFWNT9L_8tZ[118] , 
        \b11_OFWNT9L_8tZ[119] , \b11_OFWNT9L_8tZ[120] , 
        \b11_OFWNT9L_8tZ[121] , \b11_OFWNT9L_8tZ[122] , 
        \b11_OFWNT9L_8tZ[123] , \b11_OFWNT9L_8tZ[124] , 
        \b11_OFWNT9L_8tZ[125] , \b11_OFWNT9L_8tZ[126] , 
        \b11_OFWNT9L_8tZ[127] , \b11_OFWNT9L_8tZ[128] , 
        \b11_OFWNT9L_8tZ[129] , \b11_OFWNT9L_8tZ[130] , 
        \b11_OFWNT9L_8tZ[131] , \b11_OFWNT9L_8tZ[132] , 
        \b11_OFWNT9L_8tZ[133] , \b11_OFWNT9L_8tZ[134] , 
        \b11_OFWNT9L_8tZ[135] , \b11_OFWNT9L_8tZ[136] , 
        \b11_OFWNT9L_8tZ[137] , \b11_OFWNT9L_8tZ[138] , 
        \b11_OFWNT9L_8tZ[139] , \b11_OFWNT9L_8tZ[140] , 
        \b11_OFWNT9L_8tZ[141] , \b11_OFWNT9L_8tZ[142] , 
        \b11_OFWNT9L_8tZ[143] , \b11_OFWNT9L_8tZ[144] , 
        \b11_OFWNT9L_8tZ[145] , \b11_OFWNT9L_8tZ[146] , 
        \b11_OFWNT9L_8tZ[147] , \b11_OFWNT9L_8tZ[148] , 
        \b11_OFWNT9L_8tZ[149] , \b11_OFWNT9L_8tZ[150] , 
        \b11_OFWNT9L_8tZ[151] , \b11_OFWNT9L_8tZ[152] , 
        \b11_OFWNT9L_8tZ[153] , \b11_OFWNT9L_8tZ[154] , 
        \b11_OFWNT9L_8tZ[155] , \b11_OFWNT9L_8tZ[156] , 
        \b11_OFWNT9L_8tZ[157] , \b11_OFWNT9L_8tZ[158] , 
        \b11_OFWNT9L_8tZ[159] , \b11_OFWNT9L_8tZ[160] , 
        \b11_OFWNT9L_8tZ[161] , \b11_OFWNT9L_8tZ[162] , 
        \b11_OFWNT9L_8tZ[163] , \b11_OFWNT9L_8tZ[164] , 
        \b11_OFWNT9L_8tZ[165] , \b11_OFWNT9L_8tZ[166] , 
        \b11_OFWNT9L_8tZ[167] , \b11_OFWNT9L_8tZ[168] , 
        \b11_OFWNT9L_8tZ[169] , \b11_OFWNT9L_8tZ[170] , 
        \b11_OFWNT9L_8tZ[171] , \b11_OFWNT9L_8tZ[172] , 
        \b11_OFWNT9L_8tZ[173] , \b11_OFWNT9L_8tZ[174] , 
        \b11_OFWNT9L_8tZ[175] , \b11_OFWNT9L_8tZ[176] , 
        \b11_OFWNT9L_8tZ[177] , \b11_OFWNT9L_8tZ[178] , 
        \b11_OFWNT9L_8tZ[179] , \b11_OFWNT9L_8tZ[180] , 
        \b11_OFWNT9L_8tZ[181] , \b11_OFWNT9L_8tZ[182] , 
        \b11_OFWNT9L_8tZ[183] , \b11_OFWNT9L_8tZ[184] , 
        \b11_OFWNT9L_8tZ[185] , \b11_OFWNT9L_8tZ[186] , 
        \b11_OFWNT9L_8tZ[187] , \b11_OFWNT9L_8tZ[188] , 
        \b11_OFWNT9L_8tZ[189] , \b11_OFWNT9L_8tZ[190] , 
        \b11_OFWNT9L_8tZ[191] , \b11_OFWNT9L_8tZ[192] , 
        \b11_OFWNT9L_8tZ[193] , \b11_OFWNT9L_8tZ[194] , 
        \b11_OFWNT9L_8tZ[195] , \b11_OFWNT9L_8tZ[196] , 
        \b11_OFWNT9L_8tZ[197] , \b11_OFWNT9L_8tZ[198] , 
        \b11_OFWNT9L_8tZ[199] , \b11_OFWNT9L_8tZ[200] , 
        \b11_OFWNT9L_8tZ[201] , \b11_OFWNT9L_8tZ[202] , 
        \b11_OFWNT9L_8tZ[203] , \b11_OFWNT9L_8tZ[204] , 
        \b11_OFWNT9L_8tZ[205] , \b11_OFWNT9L_8tZ[206] , 
        \b11_OFWNT9L_8tZ[207] , \b11_OFWNT9L_8tZ[208] , 
        \b11_OFWNT9L_8tZ[209] , \b11_OFWNT9L_8tZ[210] , 
        \b11_OFWNT9L_8tZ[211] , \b11_OFWNT9L_8tZ[212] , 
        \b11_OFWNT9L_8tZ[213] , \b11_OFWNT9L_8tZ[214] , 
        \b11_OFWNT9L_8tZ[215] , \b11_OFWNT9L_8tZ[216] , 
        \b11_OFWNT9L_8tZ[217] , \b11_OFWNT9L_8tZ[218] , 
        \b11_OFWNT9L_8tZ[219] , \b11_OFWNT9L_8tZ[220] , 
        \b11_OFWNT9L_8tZ[221] , \b11_OFWNT9L_8tZ[222] , 
        \b11_OFWNT9L_8tZ[223] , \b11_OFWNT9L_8tZ[224] , 
        \b11_OFWNT9L_8tZ[225] , \b11_OFWNT9L_8tZ[226] , 
        \b11_OFWNT9L_8tZ[227] , \b11_OFWNT9L_8tZ[228] , 
        \b11_OFWNT9L_8tZ[229] , \b11_OFWNT9L_8tZ[230] , 
        \b11_OFWNT9L_8tZ[231] , \b11_OFWNT9L_8tZ[232] , 
        \b11_OFWNT9L_8tZ[233] , \b11_OFWNT9L_8tZ[234] , 
        \b11_OFWNT9L_8tZ[235] , \b11_OFWNT9L_8tZ[236] , 
        \b11_OFWNT9L_8tZ[237] , \b11_OFWNT9L_8tZ[238] , 
        \b11_OFWNT9L_8tZ[239] , \b11_OFWNT9L_8tZ[240] , 
        \b11_OFWNT9L_8tZ[241] , \b11_OFWNT9L_8tZ[242] , 
        \b11_OFWNT9L_8tZ[243] , \b11_OFWNT9L_8tZ[244] , 
        \b11_OFWNT9L_8tZ[245] , \b11_OFWNT9L_8tZ[246] , 
        \b11_OFWNT9L_8tZ[247] , \b11_OFWNT9L_8tZ[248] , 
        \b11_OFWNT9L_8tZ[249] , \b11_OFWNT9L_8tZ[250] , 
        \b11_OFWNT9L_8tZ[251] , \b11_OFWNT9L_8tZ[252] , 
        \b11_OFWNT9L_8tZ[253] , \b11_OFWNT9L_8tZ[254] , 
        \b11_OFWNT9L_8tZ[255] , \b11_OFWNT9L_8tZ[256] , 
        \b11_OFWNT9L_8tZ[257] , \b11_OFWNT9L_8tZ[258] , 
        \b11_OFWNT9L_8tZ[259] , \b11_OFWNT9L_8tZ[260] , 
        \b11_OFWNT9L_8tZ[261] , \b11_OFWNT9L_8tZ[262] , 
        \b11_OFWNT9L_8tZ[263] , \b11_OFWNT9L_8tZ[264] , 
        \b11_OFWNT9L_8tZ[265] , \b11_OFWNT9L_8tZ[266] , 
        \b11_OFWNT9L_8tZ[267] , \b11_OFWNT9L_8tZ[268] , 
        \b11_OFWNT9L_8tZ[269] , \b11_OFWNT9L_8tZ[270] , 
        \b11_OFWNT9L_8tZ[271] , \b11_OFWNT9L_8tZ[272] , 
        \b11_OFWNT9L_8tZ[273] , \b11_OFWNT9L_8tZ[274] , 
        \b11_OFWNT9L_8tZ[275] , \b11_OFWNT9L_8tZ[276] , 
        \b11_OFWNT9L_8tZ[277] , \b11_OFWNT9L_8tZ[278] , 
        \b11_OFWNT9L_8tZ[279] , \b11_OFWNT9L_8tZ[280] , 
        \b11_OFWNT9L_8tZ[281] , \b11_OFWNT9L_8tZ[282] , 
        \b11_OFWNT9L_8tZ[283] , \b11_OFWNT9L_8tZ[284] , 
        \b11_OFWNT9L_8tZ[285] , \b11_OFWNT9L_8tZ[286] , 
        \b11_OFWNT9L_8tZ[287] , \b11_OFWNT9L_8tZ[288] , 
        \b11_OFWNT9L_8tZ[289] , \b11_OFWNT9L_8tZ[290] , 
        \b11_OFWNT9L_8tZ[291] , \b11_OFWNT9L_8tZ[292] , 
        \b11_OFWNT9L_8tZ[293] , \b11_OFWNT9L_8tZ[294] , 
        \b11_OFWNT9L_8tZ[295] , \b11_OFWNT9L_8tZ[296] , 
        \b11_OFWNT9L_8tZ[297] , \b11_OFWNT9L_8tZ[298] , 
        \b11_OFWNT9L_8tZ[299] , \b11_OFWNT9L_8tZ[300] , 
        \b11_OFWNT9L_8tZ[301] , \b11_OFWNT9L_8tZ[302] , 
        \b11_OFWNT9L_8tZ[303] , \b11_OFWNT9L_8tZ[304] , 
        \b11_OFWNT9L_8tZ[305] , \b11_OFWNT9L_8tZ[306] , 
        \b11_OFWNT9L_8tZ[307] , \b11_OFWNT9L_8tZ[308] , 
        \b11_OFWNT9L_8tZ[309] , \b11_OFWNT9L_8tZ[310] , 
        \b11_OFWNT9L_8tZ[311] , \b11_OFWNT9L_8tZ[312] , 
        \b11_OFWNT9L_8tZ[313] , \b11_OFWNT9L_8tZ[314] , 
        \b11_OFWNT9L_8tZ[315] , \b11_OFWNT9L_8tZ[316] , 
        \b11_OFWNT9L_8tZ[317] , \b11_OFWNT9L_8tZ[318] , 
        \b11_OFWNT9L_8tZ[319] , \b11_OFWNT9L_8tZ[320] , 
        \b11_OFWNT9L_8tZ[321] , \b11_OFWNT9L_8tZ[322] , 
        \b11_OFWNT9L_8tZ[323] , \b11_OFWNT9L_8tZ[324] , 
        \b11_OFWNT9L_8tZ[325] , \b11_OFWNT9L_8tZ[326] , 
        \b11_OFWNT9L_8tZ[327] , \b11_OFWNT9L_8tZ[328] , 
        \b11_OFWNT9L_8tZ[329] , \b11_OFWNT9L_8tZ[330] , 
        \b11_OFWNT9L_8tZ[331] , \b11_OFWNT9L_8tZ[332] , 
        \b11_OFWNT9L_8tZ[333] , \b11_OFWNT9L_8tZ[334] , 
        \b11_OFWNT9L_8tZ[335] , \b11_OFWNT9L_8tZ[336] , 
        \b11_OFWNT9L_8tZ[337] , \b11_OFWNT9L_8tZ[338] , 
        \b11_OFWNT9L_8tZ[339] , \b11_OFWNT9L_8tZ[340] , 
        \b11_OFWNT9L_8tZ[341] , \b11_OFWNT9L_8tZ[342] , 
        \b11_OFWNT9L_8tZ[343] , \b11_OFWNT9L_8tZ[344] , 
        \b11_OFWNT9L_8tZ[345] , \b11_OFWNT9L_8tZ[346] , 
        \b11_OFWNT9L_8tZ[347] , \b11_OFWNT9L_8tZ[348] , 
        \b11_OFWNT9L_8tZ[349] , \b11_OFWNT9L_8tZ[350] , 
        \b11_OFWNT9L_8tZ[351] , \b11_OFWNT9L_8tZ[352] , 
        \b11_OFWNT9L_8tZ[353] , \b11_OFWNT9L_8tZ[354] , 
        \b11_OFWNT9L_8tZ[355] , \b11_OFWNT9L_8tZ[356] , 
        \b11_OFWNT9L_8tZ[357] , \b11_OFWNT9L_8tZ[358] , 
        \b11_OFWNT9L_8tZ[359] , \b11_OFWNT9L_8tZ[360] , 
        \b11_OFWNT9L_8tZ[361] , \b11_OFWNT9L_8tZ[362] , 
        \b11_OFWNT9L_8tZ[363] , \b11_OFWNT9L_8tZ[364] , 
        \b11_OFWNT9L_8tZ[365] , \b11_OFWNT9L_8tZ[366] , 
        \b11_OFWNT9L_8tZ[367] , \b11_OFWNT9L_8tZ[368] , 
        \b11_OFWNT9L_8tZ[369] , \b11_OFWNT9L_8tZ[370] , 
        \b11_OFWNT9L_8tZ[371] , \b11_OFWNT9L_8tZ[372] , 
        \b11_OFWNT9L_8tZ[373] , \b11_OFWNT9L_8tZ[374] , 
        \b11_OFWNT9L_8tZ[375] , \b11_OFWNT9L_8tZ[376] , b8_SoWGfWYY, 
        b8_SoWGfWYY_i, b11_PSyil9s_FMZ;
    
    SLE \mdiclink_reg[291]  (.D(temp3[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[291]_net_1 ));
    SLE \mdiclink_reg[279]  (.D(temp2[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[279]_net_1 ));
    SLE \mdiclink_reg[162]  (.D(dds_cos[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[162]_net_1 ));
    SLE \mdiclink_reg[346]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[346]_net_1 ));
    SLE \mdiclink_reg[89]  (.D(\data_from_adc[5] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[89]_net_1 ));
    SLE \mdiclink_reg[117]  (.D(\data_from_adc[3] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[117]_net_1 ));
    SLE \mdiclink_reg[184]  (.D(fpga_count[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[184]_net_1 ));
    SLE \mdiclink_reg[116]  (.D(\data_from_adc[3] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[116]_net_1 ));
    SLE \mdiclink_reg[110]  (.D(\data_from_adc[3] [11]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[110]_net_1 ));
    SLE \mdiclink_reg[171]  (.D(dds_sin[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[171]_net_1 ));
    SLE \mdiclink_reg[90]  (.D(\data_from_adc[5] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[90]_net_1 ));
    SLE \mdiclink_reg[366]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[366]_net_1 ));
    SLE \mdiclink_reg[327]  (.D(temp_count[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[327]_net_1 ));
    SLE \mdiclink_reg[319]  (.D(temp_count[18]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[319]_net_1 ));
    SLE \mdiclink_reg[97]  (.D(\data_from_adc[5] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[97]_net_1 ));
    SLE \mdiclink_reg[240]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[240]_net_1 ));
    SLE \mdiclink_reg[108]  (.D(\data_from_adc[4] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[108]_net_1 ));
    SLE \mdiclink_reg[216]  (.D(fr_adc_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[216]_net_1 ));
    SLE \mdiclink_reg[155]  (.D(\data_from_adc[0] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[155]_net_1 ));
    SLE \mdiclink_reg[134]  (.D(\data_from_adc[1] [11]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[134]_net_1 ));
    SLE \mdiclink_reg[281]  (.D(temp2[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[281]_net_1 ));
    SLE \mdiclink_reg[208]  (.D(fr_adc_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[208]_net_1 ));
    SLE \mdiclink_reg[335]  (.D(temp_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[335]_net_1 ));
    SLE \mdiclink_reg[204]  (.D(fpga_shift_2[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[204]_net_1 ));
    SLE \mdiclink_reg[61]  (.D(\data_from_adc[8] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[61]_net_1 ));
    SLE \mdiclink_reg[129]  (.D(\data_from_adc[2] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[129]_net_1 ));
    SLE \mdiclink_reg[260]  (.D(temp1[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[260]_net_1 ));
    SLE \mdiclink_reg[310]  (.D(temp_count[27]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[310]_net_1 ));
    SLE \mdiclink_reg[231]  (.D(freq_14), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[231]_net_1 ));
    SLE \mdiclink_reg[203]  (.D(fpga_shift_2[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[203]_net_1 ));
    SLE \mdiclink_reg[172]  (.D(dds_sin[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[172]_net_1 ));
    SLE \mdiclink_reg[2]  (.D(BW_c[12]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[2]_net_1 ));
    SLE \mdiclink_reg[85]  (.D(\data_from_adc[6] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[85]_net_1 ));
    SLE \mdiclink_reg[292]  (.D(temp3[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[292]_net_1 ));
    SLE \mdiclink_reg[49]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[49]_net_1 ));
    SLE \mdiclink_reg[245]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[245]_net_1 ));
    SLE \mdiclink_reg[331]  (.D(temp_count[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[331]_net_1 ));
    SLE \mdiclink_reg[304]  (.D(temp3[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[304]_net_1 ));
    SLE \mdiclink_reg[376]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[376]_net_1 ));
    SLE \mdiclink_reg[127]  (.D(\data_from_adc[2] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[127]_net_1 ));
    SLE \mdiclink_reg[63]  (.D(\data_from_adc[7] [10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[63]_net_1 ));
    SLE \mdiclink_reg[357]  (.D(VCC_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[357]_net_1 ));
    SLE \mdiclink_reg[297]  (.D(temp3[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[297]_net_1 ));
    SLE \mdiclink_reg[126]  (.D(\data_from_adc[2] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[126]_net_1 ));
    SLE \mdiclink_reg[120]  (.D(\data_from_adc[3] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[120]_net_1 ));
    SLE \mdiclink_reg[265]  (.D(temp1[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[265]_net_1 ));
    SLE \mdiclink_reg[80]  (.D(\data_from_adc[6] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[80]_net_1 ));
    SLE \mdiclink_reg[329]  (.D(temp_count[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[329]_net_1 ));
    SLE \mdiclink_reg[270]  (.D(temp1[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[270]_net_1 ));
    SLE \mdiclink_reg[159]  (.D(dds_cos[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[159]_net_1 ));
    SLE \mdiclink_reg[52]  (.D(\data_from_adc[8] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[52]_net_1 ));
    SLE \mdiclink_reg[226]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[226]_net_1 ));
    SLE \mdiclink_reg[87]  (.D(\data_from_adc[5] [10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[87]_net_1 ));
    SLE \mdiclink_reg[313]  (.D(temp_count[24]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[313]_net_1 ));
    SLE \mdiclink_reg[68]  (.D(\data_from_adc[7] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[68]_net_1 ));
    SLE \mdiclink_reg[31]  (.D(clk_dac2), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[31]_net_1 ));
    SLE \mdiclink_reg[282]  (.D(temp2[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[282]_net_1 ));
    SLE \mdiclink_reg[103]  (.D(\data_from_adc[4] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[103]_net_1 ));
    SLE \mdiclink_reg[332]  (.D(temp_count[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[332]_net_1 ));
    SLE \mdiclink_reg[320]  (.D(temp_count[17]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[320]_net_1 ));
    SLE \mdiclink_reg[66]  (.D(\data_from_adc[7] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[66]_net_1 ));
    SLE \mdiclink_reg[45]  (.D(dac_count[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[45]_net_1 ));
    SLE \mdiclink_reg[287]  (.D(temp2[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[287]_net_1 ));
    SLE \mdiclink_reg[232]  (.D(freq_13), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[232]_net_1 ));
    SLE \mdiclink_reg[157]  (.D(\data_from_adc[0] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[157]_net_1 ));
    SLE \mdiclink_reg[54]  (.D(\data_from_adc[8] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[54]_net_1 ));
    SLE \mdiclink_reg[156]  (.D(\data_from_adc[0] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[156]_net_1 ));
    SLE \mdiclink_reg[275]  (.D(temp2[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[275]_net_1 ));
    SLE \mdiclink_reg[150]  (.D(\data_from_adc[0] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[150]_net_1 ));
    SLE \mdiclink_reg[237]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[237]_net_1 ));
    SLE \mdiclink_reg[33]  (.D(dac1_db_c[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[33]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \mdiclink_reg[40]  (.D(dac1_db_c[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[40]_net_1 ));
    SLE \mdiclink_reg[359]  (.D(freq_10), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[359]_net_1 ));
    SLE \mdiclink_reg[105]  (.D(\data_from_adc[4] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[105]_net_1 ));
    SLE \mdiclink_reg[256]  (.D(temp1[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[256]_net_1 ));
    SLE \mdiclink_reg[47]  (.D(dac_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[47]_net_1 ));
    SLE \mdiclink_reg[299]  (.D(temp3[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[299]_net_1 ));
    SLE \mdiclink_reg[148]  (.D(\data_from_adc[0] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[148]_net_1 ));
    SLE \mdiclink_reg[248]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[248]_net_1 ));
    SLE \mdiclink_reg[114]  (.D(\data_from_adc[3] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[114]_net_1 ));
    SLE \mdiclink_reg[244]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[244]_net_1 ));
    SLE \mdiclink_reg[350]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[350]_net_1 ));
    SLE \mdiclink_reg[323]  (.D(temp_count[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[323]_net_1 ));
    SLE \mdiclink_reg[38]  (.D(dac1_db_c[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[38]_net_1 ));
    SLE \mdiclink_reg[315]  (.D(temp_count[22]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[315]_net_1 ));
    SLE \mdiclink_reg[168]  (.D(dds_sin[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[168]_net_1 ));
    SLE \mdiclink_reg[191]  (.D(fpga_shift_2[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[191]_net_1 ));
    SLE \mdiclink_reg[268]  (.D(temp1[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[268]_net_1 ));
    SLE \mdiclink_reg[264]  (.D(temp1[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[264]_net_1 ));
    SLE \mdiclink_reg[36]  (.D(dac1_db_c[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[36]_net_1 ));
    SLE \mdiclink_reg[243]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[243]_net_1 ));
    SLE \mdiclink_reg[21]  (.D(BW_out_c[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[21]_net_1 ));
    SLE \mdiclink_reg[211]  (.D(fr_adc_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[211]_net_1 ));
    b3_12m_x_0 b8_12m_IFLY (.b6_Ocm0rW_0_0_o2({\b6_Ocm0rW_0_0_o2[2] }), 
        .b13_nAzGfFM_sLsv3({\b13_nAzGfFM_sLsv3[1] }), .IICE_comm2iice({
        IICE_comm2iice[11], IICE_comm2iice[10], IICE_comm2iice[9], 
        IICE_comm2iice[8]}), .mdiclink_reg({\mdiclink_reg[376]_net_1 , 
        \mdiclink_reg[375]_net_1 , \mdiclink_reg[374]_net_1 , 
        \mdiclink_reg[373]_net_1 , \mdiclink_reg[372]_net_1 , 
        \mdiclink_reg[371]_net_1 , \mdiclink_reg[370]_net_1 , 
        \mdiclink_reg[369]_net_1 , \mdiclink_reg[368]_net_1 , 
        \mdiclink_reg[367]_net_1 , \mdiclink_reg[366]_net_1 , 
        \mdiclink_reg[365]_net_1 , \mdiclink_reg[364]_net_1 , 
        \mdiclink_reg[363]_net_1 , \mdiclink_reg[362]_net_1 , 
        \mdiclink_reg[361]_net_1 , \mdiclink_reg[360]_net_1 , 
        \mdiclink_reg[359]_net_1 , \mdiclink_reg[358]_net_1 , 
        \mdiclink_reg[357]_net_1 , \mdiclink_reg[356]_net_1 , 
        \mdiclink_reg[355]_net_1 , \mdiclink_reg[354]_net_1 , 
        \mdiclink_reg[353]_net_1 , \mdiclink_reg[352]_net_1 , 
        \mdiclink_reg[351]_net_1 , \mdiclink_reg[350]_net_1 , 
        \mdiclink_reg[349]_net_1 , \mdiclink_reg[348]_net_1 , 
        \mdiclink_reg[347]_net_1 , \mdiclink_reg[346]_net_1 , 
        \mdiclink_reg[345]_net_1 , \mdiclink_reg[344]_net_1 , 
        \mdiclink_reg[343]_net_1 , \mdiclink_reg[342]_net_1 , 
        \mdiclink_reg[341]_net_1 , \mdiclink_reg[340]_net_1 , 
        \mdiclink_reg[339]_net_1 , \mdiclink_reg[338]_net_1 , 
        \mdiclink_reg[337]_net_1 , \mdiclink_reg[336]_net_1 , 
        \mdiclink_reg[335]_net_1 , \mdiclink_reg[334]_net_1 , 
        \mdiclink_reg[333]_net_1 , \mdiclink_reg[332]_net_1 , 
        \mdiclink_reg[331]_net_1 , \mdiclink_reg[330]_net_1 , 
        \mdiclink_reg[329]_net_1 , \mdiclink_reg[328]_net_1 , 
        \mdiclink_reg[327]_net_1 , \mdiclink_reg[326]_net_1 , 
        \mdiclink_reg[325]_net_1 , \mdiclink_reg[324]_net_1 , 
        \mdiclink_reg[323]_net_1 , \mdiclink_reg[322]_net_1 , 
        \mdiclink_reg[321]_net_1 , \mdiclink_reg[320]_net_1 , 
        \mdiclink_reg[319]_net_1 , \mdiclink_reg[318]_net_1 , 
        \mdiclink_reg[317]_net_1 , \mdiclink_reg[316]_net_1 , 
        \mdiclink_reg[315]_net_1 , \mdiclink_reg[314]_net_1 , 
        \mdiclink_reg[313]_net_1 , \mdiclink_reg[312]_net_1 , 
        \mdiclink_reg[311]_net_1 , \mdiclink_reg[310]_net_1 , 
        \mdiclink_reg[309]_net_1 , \mdiclink_reg[308]_net_1 , 
        \mdiclink_reg[307]_net_1 , \mdiclink_reg[306]_net_1 , 
        \mdiclink_reg[305]_net_1 , \mdiclink_reg[304]_net_1 , 
        \mdiclink_reg[303]_net_1 , \mdiclink_reg[302]_net_1 , 
        \mdiclink_reg[301]_net_1 , \mdiclink_reg[300]_net_1 , 
        \mdiclink_reg[299]_net_1 , \mdiclink_reg[298]_net_1 , 
        \mdiclink_reg[297]_net_1 , \mdiclink_reg[296]_net_1 , 
        \mdiclink_reg[295]_net_1 , \mdiclink_reg[294]_net_1 , 
        \mdiclink_reg[293]_net_1 , \mdiclink_reg[292]_net_1 , 
        \mdiclink_reg[291]_net_1 , \mdiclink_reg[290]_net_1 , 
        \mdiclink_reg[289]_net_1 , \mdiclink_reg[288]_net_1 , 
        \mdiclink_reg[287]_net_1 , \mdiclink_reg[286]_net_1 , 
        \mdiclink_reg[285]_net_1 , \mdiclink_reg[284]_net_1 , 
        \mdiclink_reg[283]_net_1 , \mdiclink_reg[282]_net_1 , 
        \mdiclink_reg[281]_net_1 , \mdiclink_reg[280]_net_1 , 
        \mdiclink_reg[279]_net_1 , \mdiclink_reg[278]_net_1 , 
        \mdiclink_reg[277]_net_1 , \mdiclink_reg[276]_net_1 , 
        \mdiclink_reg[275]_net_1 , \mdiclink_reg[274]_net_1 , 
        \mdiclink_reg[273]_net_1 , \mdiclink_reg[272]_net_1 , 
        \mdiclink_reg[271]_net_1 , \mdiclink_reg[270]_net_1 , 
        \mdiclink_reg[269]_net_1 , \mdiclink_reg[268]_net_1 , 
        \mdiclink_reg[267]_net_1 , \mdiclink_reg[266]_net_1 , 
        \mdiclink_reg[265]_net_1 , \mdiclink_reg[264]_net_1 , 
        \mdiclink_reg[263]_net_1 , \mdiclink_reg[262]_net_1 , 
        \mdiclink_reg[261]_net_1 , \mdiclink_reg[260]_net_1 , 
        \mdiclink_reg[259]_net_1 , \mdiclink_reg[258]_net_1 , 
        \mdiclink_reg[257]_net_1 , \mdiclink_reg[256]_net_1 , 
        \mdiclink_reg[255]_net_1 , \mdiclink_reg[254]_net_1 , 
        \mdiclink_reg[253]_net_1 , \mdiclink_reg[252]_net_1 , 
        \mdiclink_reg[251]_net_1 , \mdiclink_reg[250]_net_1 , 
        \mdiclink_reg[249]_net_1 , \mdiclink_reg[248]_net_1 , 
        \mdiclink_reg[247]_net_1 , \mdiclink_reg[246]_net_1 , 
        \mdiclink_reg[245]_net_1 , \mdiclink_reg[244]_net_1 , 
        \mdiclink_reg[243]_net_1 , \mdiclink_reg[242]_net_1 , 
        \mdiclink_reg[241]_net_1 , \mdiclink_reg[240]_net_1 , 
        \mdiclink_reg[239]_net_1 , \mdiclink_reg[238]_net_1 , 
        \mdiclink_reg[237]_net_1 , \mdiclink_reg[236]_net_1 , 
        \mdiclink_reg[235]_net_1 , \mdiclink_reg[234]_net_1 , 
        \mdiclink_reg[233]_net_1 , \mdiclink_reg[232]_net_1 , 
        \mdiclink_reg[231]_net_1 , \mdiclink_reg[230]_net_1 , 
        \mdiclink_reg[229]_net_1 , \mdiclink_reg[228]_net_1 , 
        \mdiclink_reg[227]_net_1 , \mdiclink_reg[226]_net_1 , 
        \mdiclink_reg[225]_net_1 , \mdiclink_reg[224]_net_1 , 
        \mdiclink_reg[223]_net_1 , \mdiclink_reg[222]_net_1 , 
        \mdiclink_reg[221]_net_1 , \mdiclink_reg[220]_net_1 , 
        \mdiclink_reg[219]_net_1 , \mdiclink_reg[218]_net_1 , 
        \mdiclink_reg[217]_net_1 , \mdiclink_reg[216]_net_1 , 
        \mdiclink_reg[215]_net_1 , \mdiclink_reg[214]_net_1 , 
        \mdiclink_reg[213]_net_1 , \mdiclink_reg[212]_net_1 , 
        \mdiclink_reg[211]_net_1 , \mdiclink_reg[210]_net_1 , 
        \mdiclink_reg[209]_net_1 , \mdiclink_reg[208]_net_1 , 
        \mdiclink_reg[207]_net_1 , \mdiclink_reg[206]_net_1 , 
        \mdiclink_reg[205]_net_1 , \mdiclink_reg[204]_net_1 , 
        \mdiclink_reg[203]_net_1 , \mdiclink_reg[202]_net_1 , 
        \mdiclink_reg[201]_net_1 , \mdiclink_reg[200]_net_1 , 
        \mdiclink_reg[199]_net_1 , \mdiclink_reg[198]_net_1 , 
        \mdiclink_reg[197]_net_1 , \mdiclink_reg[196]_net_1 , 
        \mdiclink_reg[195]_net_1 , \mdiclink_reg[194]_net_1 , 
        \mdiclink_reg[193]_net_1 , \mdiclink_reg[192]_net_1 , 
        \mdiclink_reg[191]_net_1 , \mdiclink_reg[190]_net_1 , 
        \mdiclink_reg[189]_net_1 , \mdiclink_reg[188]_net_1 , 
        \mdiclink_reg[187]_net_1 , \mdiclink_reg[186]_net_1 , 
        \mdiclink_reg[185]_net_1 , \mdiclink_reg[184]_net_1 , 
        \mdiclink_reg[183]_net_1 , \mdiclink_reg[182]_net_1 , 
        \mdiclink_reg[181]_net_1 , \mdiclink_reg[180]_net_1 , 
        \mdiclink_reg[179]_net_1 , \mdiclink_reg[178]_net_1 , 
        \mdiclink_reg[177]_net_1 , \mdiclink_reg[176]_net_1 , 
        \mdiclink_reg[175]_net_1 , \mdiclink_reg[174]_net_1 , 
        \mdiclink_reg[173]_net_1 , \mdiclink_reg[172]_net_1 , 
        \mdiclink_reg[171]_net_1 , \mdiclink_reg[170]_net_1 , 
        \mdiclink_reg[169]_net_1 , \mdiclink_reg[168]_net_1 , 
        \mdiclink_reg[167]_net_1 , \mdiclink_reg[166]_net_1 , 
        \mdiclink_reg[165]_net_1 , \mdiclink_reg[164]_net_1 , 
        \mdiclink_reg[163]_net_1 , \mdiclink_reg[162]_net_1 , 
        \mdiclink_reg[161]_net_1 , \mdiclink_reg[160]_net_1 , 
        \mdiclink_reg[159]_net_1 , \mdiclink_reg[158]_net_1 , 
        \mdiclink_reg[157]_net_1 , \mdiclink_reg[156]_net_1 , 
        \mdiclink_reg[155]_net_1 , \mdiclink_reg[154]_net_1 , 
        \mdiclink_reg[153]_net_1 , \mdiclink_reg[152]_net_1 , 
        \mdiclink_reg[151]_net_1 , \mdiclink_reg[150]_net_1 , 
        \mdiclink_reg[149]_net_1 , \mdiclink_reg[148]_net_1 , 
        \mdiclink_reg[147]_net_1 , \mdiclink_reg[146]_net_1 , 
        \mdiclink_reg[145]_net_1 , \mdiclink_reg[144]_net_1 , 
        \mdiclink_reg[143]_net_1 , \mdiclink_reg[142]_net_1 , 
        \mdiclink_reg[141]_net_1 , \mdiclink_reg[140]_net_1 , 
        \mdiclink_reg[139]_net_1 , \mdiclink_reg[138]_net_1 , 
        \mdiclink_reg[137]_net_1 , \mdiclink_reg[136]_net_1 , 
        \mdiclink_reg[135]_net_1 , \mdiclink_reg[134]_net_1 , 
        \mdiclink_reg[133]_net_1 , \mdiclink_reg[132]_net_1 , 
        \mdiclink_reg[131]_net_1 , \mdiclink_reg[130]_net_1 , 
        \mdiclink_reg[129]_net_1 , \mdiclink_reg[128]_net_1 , 
        \mdiclink_reg[127]_net_1 , \mdiclink_reg[126]_net_1 , 
        \mdiclink_reg[125]_net_1 , \mdiclink_reg[124]_net_1 , 
        \mdiclink_reg[123]_net_1 , \mdiclink_reg[122]_net_1 , 
        \mdiclink_reg[121]_net_1 , \mdiclink_reg[120]_net_1 , 
        \mdiclink_reg[119]_net_1 , \mdiclink_reg[118]_net_1 , 
        \mdiclink_reg[117]_net_1 , \mdiclink_reg[116]_net_1 , 
        \mdiclink_reg[115]_net_1 , \mdiclink_reg[114]_net_1 , 
        \mdiclink_reg[113]_net_1 , \mdiclink_reg[112]_net_1 , 
        \mdiclink_reg[111]_net_1 , \mdiclink_reg[110]_net_1 , 
        \mdiclink_reg[109]_net_1 , \mdiclink_reg[108]_net_1 , 
        \mdiclink_reg[107]_net_1 , \mdiclink_reg[106]_net_1 , 
        \mdiclink_reg[105]_net_1 , \mdiclink_reg[104]_net_1 , 
        \mdiclink_reg[103]_net_1 , \mdiclink_reg[102]_net_1 , 
        \mdiclink_reg[101]_net_1 , \mdiclink_reg[100]_net_1 , 
        \mdiclink_reg[99]_net_1 , \mdiclink_reg[98]_net_1 , 
        \mdiclink_reg[97]_net_1 , \mdiclink_reg[96]_net_1 , 
        \mdiclink_reg[95]_net_1 , \mdiclink_reg[94]_net_1 , 
        \mdiclink_reg[93]_net_1 , \mdiclink_reg[92]_net_1 , 
        \mdiclink_reg[91]_net_1 , \mdiclink_reg[90]_net_1 , 
        \mdiclink_reg[89]_net_1 , \mdiclink_reg[88]_net_1 , 
        \mdiclink_reg[87]_net_1 , \mdiclink_reg[86]_net_1 , 
        \mdiclink_reg[85]_net_1 , \mdiclink_reg[84]_net_1 , 
        \mdiclink_reg[83]_net_1 , \mdiclink_reg[82]_net_1 , 
        \mdiclink_reg[81]_net_1 , \mdiclink_reg[80]_net_1 , 
        \mdiclink_reg[79]_net_1 , \mdiclink_reg[78]_net_1 , 
        \mdiclink_reg[77]_net_1 , \mdiclink_reg[76]_net_1 , 
        \mdiclink_reg[75]_net_1 , \mdiclink_reg[74]_net_1 , 
        \mdiclink_reg[73]_net_1 , \mdiclink_reg[72]_net_1 , 
        \mdiclink_reg[71]_net_1 , \mdiclink_reg[70]_net_1 , 
        \mdiclink_reg[69]_net_1 , \mdiclink_reg[68]_net_1 , 
        \mdiclink_reg[67]_net_1 , \mdiclink_reg[66]_net_1 , 
        \mdiclink_reg[65]_net_1 , \mdiclink_reg[64]_net_1 , 
        \mdiclink_reg[63]_net_1 , \mdiclink_reg[62]_net_1 , 
        \mdiclink_reg[61]_net_1 , \mdiclink_reg[60]_net_1 , 
        \mdiclink_reg[59]_net_1 , \mdiclink_reg[58]_net_1 , 
        \mdiclink_reg[57]_net_1 , \mdiclink_reg[56]_net_1 , 
        \mdiclink_reg[55]_net_1 , \mdiclink_reg[54]_net_1 , 
        \mdiclink_reg[53]_net_1 , \mdiclink_reg[52]_net_1 , 
        \mdiclink_reg[51]_net_1 , \mdiclink_reg[50]_net_1 , 
        \mdiclink_reg[49]_net_1 , \mdiclink_reg[48]_net_1 , 
        \mdiclink_reg[47]_net_1 , \mdiclink_reg[46]_net_1 , 
        \mdiclink_reg[45]_net_1 , \mdiclink_reg[44]_net_1 , 
        \mdiclink_reg[43]_net_1 , \mdiclink_reg[42]_net_1 , 
        \mdiclink_reg[41]_net_1 , \mdiclink_reg[40]_net_1 , 
        \mdiclink_reg[39]_net_1 , \mdiclink_reg[38]_net_1 , 
        \mdiclink_reg[37]_net_1 , \mdiclink_reg[36]_net_1 , 
        \mdiclink_reg[35]_net_1 , \mdiclink_reg[34]_net_1 , 
        \mdiclink_reg[33]_net_1 , \mdiclink_reg[32]_net_1 , 
        \mdiclink_reg[31]_net_1 , \mdiclink_reg[30]_net_1 , 
        \mdiclink_reg[29]_net_1 , \mdiclink_reg[28]_net_1 , 
        \mdiclink_reg[27]_net_1 , \mdiclink_reg[26]_net_1 , 
        \mdiclink_reg[25]_net_1 , \mdiclink_reg[24]_net_1 , 
        \mdiclink_reg[23]_net_1 , \mdiclink_reg[22]_net_1 , 
        \mdiclink_reg[21]_net_1 , \mdiclink_reg[20]_net_1 , 
        \mdiclink_reg[19]_net_1 , \mdiclink_reg[18]_net_1 , 
        \mdiclink_reg[17]_net_1 , \mdiclink_reg[16]_net_1 , 
        \mdiclink_reg[15]_net_1 , \mdiclink_reg[14]_net_1 , 
        \mdiclink_reg[13]_net_1 , \mdiclink_reg[12]_net_1 , 
        \mdiclink_reg[11]_net_1 , \mdiclink_reg[10]_net_1 , 
        \mdiclink_reg[9]_net_1 , \mdiclink_reg[8]_net_1 , 
        \mdiclink_reg[7]_net_1 , \mdiclink_reg[6]_net_1 , 
        \mdiclink_reg[5]_net_1 , \mdiclink_reg[4]_net_1 , 
        \mdiclink_reg[3]_net_1 , \mdiclink_reg[2]_net_1 , 
        \mdiclink_reg[1]_net_1 , \mdiclink_reg[0]_net_1 }), 
        .b11_OFWNT9L_8tZ({\b11_OFWNT9L_8tZ[376] , 
        \b11_OFWNT9L_8tZ[375] , \b11_OFWNT9L_8tZ[374] , 
        \b11_OFWNT9L_8tZ[373] , \b11_OFWNT9L_8tZ[372] , 
        \b11_OFWNT9L_8tZ[371] , \b11_OFWNT9L_8tZ[370] , 
        \b11_OFWNT9L_8tZ[369] , \b11_OFWNT9L_8tZ[368] , 
        \b11_OFWNT9L_8tZ[367] , \b11_OFWNT9L_8tZ[366] , 
        \b11_OFWNT9L_8tZ[365] , \b11_OFWNT9L_8tZ[364] , 
        \b11_OFWNT9L_8tZ[363] , \b11_OFWNT9L_8tZ[362] , 
        \b11_OFWNT9L_8tZ[361] , \b11_OFWNT9L_8tZ[360] , 
        \b11_OFWNT9L_8tZ[359] , \b11_OFWNT9L_8tZ[358] , 
        \b11_OFWNT9L_8tZ[357] , \b11_OFWNT9L_8tZ[356] , 
        \b11_OFWNT9L_8tZ[355] , \b11_OFWNT9L_8tZ[354] , 
        \b11_OFWNT9L_8tZ[353] , \b11_OFWNT9L_8tZ[352] , 
        \b11_OFWNT9L_8tZ[351] , \b11_OFWNT9L_8tZ[350] , 
        \b11_OFWNT9L_8tZ[349] , \b11_OFWNT9L_8tZ[348] , 
        \b11_OFWNT9L_8tZ[347] , \b11_OFWNT9L_8tZ[346] , 
        \b11_OFWNT9L_8tZ[345] , \b11_OFWNT9L_8tZ[344] , 
        \b11_OFWNT9L_8tZ[343] , \b11_OFWNT9L_8tZ[342] , 
        \b11_OFWNT9L_8tZ[341] , \b11_OFWNT9L_8tZ[340] , 
        \b11_OFWNT9L_8tZ[339] , \b11_OFWNT9L_8tZ[338] , 
        \b11_OFWNT9L_8tZ[337] , \b11_OFWNT9L_8tZ[336] , 
        \b11_OFWNT9L_8tZ[335] , \b11_OFWNT9L_8tZ[334] , 
        \b11_OFWNT9L_8tZ[333] , \b11_OFWNT9L_8tZ[332] , 
        \b11_OFWNT9L_8tZ[331] , \b11_OFWNT9L_8tZ[330] , 
        \b11_OFWNT9L_8tZ[329] , \b11_OFWNT9L_8tZ[328] , 
        \b11_OFWNT9L_8tZ[327] , \b11_OFWNT9L_8tZ[326] , 
        \b11_OFWNT9L_8tZ[325] , \b11_OFWNT9L_8tZ[324] , 
        \b11_OFWNT9L_8tZ[323] , \b11_OFWNT9L_8tZ[322] , 
        \b11_OFWNT9L_8tZ[321] , \b11_OFWNT9L_8tZ[320] , 
        \b11_OFWNT9L_8tZ[319] , \b11_OFWNT9L_8tZ[318] , 
        \b11_OFWNT9L_8tZ[317] , \b11_OFWNT9L_8tZ[316] , 
        \b11_OFWNT9L_8tZ[315] , \b11_OFWNT9L_8tZ[314] , 
        \b11_OFWNT9L_8tZ[313] , \b11_OFWNT9L_8tZ[312] , 
        \b11_OFWNT9L_8tZ[311] , \b11_OFWNT9L_8tZ[310] , 
        \b11_OFWNT9L_8tZ[309] , \b11_OFWNT9L_8tZ[308] , 
        \b11_OFWNT9L_8tZ[307] , \b11_OFWNT9L_8tZ[306] , 
        \b11_OFWNT9L_8tZ[305] , \b11_OFWNT9L_8tZ[304] , 
        \b11_OFWNT9L_8tZ[303] , \b11_OFWNT9L_8tZ[302] , 
        \b11_OFWNT9L_8tZ[301] , \b11_OFWNT9L_8tZ[300] , 
        \b11_OFWNT9L_8tZ[299] , \b11_OFWNT9L_8tZ[298] , 
        \b11_OFWNT9L_8tZ[297] , \b11_OFWNT9L_8tZ[296] , 
        \b11_OFWNT9L_8tZ[295] , \b11_OFWNT9L_8tZ[294] , 
        \b11_OFWNT9L_8tZ[293] , \b11_OFWNT9L_8tZ[292] , 
        \b11_OFWNT9L_8tZ[291] , \b11_OFWNT9L_8tZ[290] , 
        \b11_OFWNT9L_8tZ[289] , \b11_OFWNT9L_8tZ[288] , 
        \b11_OFWNT9L_8tZ[287] , \b11_OFWNT9L_8tZ[286] , 
        \b11_OFWNT9L_8tZ[285] , \b11_OFWNT9L_8tZ[284] , 
        \b11_OFWNT9L_8tZ[283] , \b11_OFWNT9L_8tZ[282] , 
        \b11_OFWNT9L_8tZ[281] , \b11_OFWNT9L_8tZ[280] , 
        \b11_OFWNT9L_8tZ[279] , \b11_OFWNT9L_8tZ[278] , 
        \b11_OFWNT9L_8tZ[277] , \b11_OFWNT9L_8tZ[276] , 
        \b11_OFWNT9L_8tZ[275] , \b11_OFWNT9L_8tZ[274] , 
        \b11_OFWNT9L_8tZ[273] , \b11_OFWNT9L_8tZ[272] , 
        \b11_OFWNT9L_8tZ[271] , \b11_OFWNT9L_8tZ[270] , 
        \b11_OFWNT9L_8tZ[269] , \b11_OFWNT9L_8tZ[268] , 
        \b11_OFWNT9L_8tZ[267] , \b11_OFWNT9L_8tZ[266] , 
        \b11_OFWNT9L_8tZ[265] , \b11_OFWNT9L_8tZ[264] , 
        \b11_OFWNT9L_8tZ[263] , \b11_OFWNT9L_8tZ[262] , 
        \b11_OFWNT9L_8tZ[261] , \b11_OFWNT9L_8tZ[260] , 
        \b11_OFWNT9L_8tZ[259] , \b11_OFWNT9L_8tZ[258] , 
        \b11_OFWNT9L_8tZ[257] , \b11_OFWNT9L_8tZ[256] , 
        \b11_OFWNT9L_8tZ[255] , \b11_OFWNT9L_8tZ[254] , 
        \b11_OFWNT9L_8tZ[253] , \b11_OFWNT9L_8tZ[252] , 
        \b11_OFWNT9L_8tZ[251] , \b11_OFWNT9L_8tZ[250] , 
        \b11_OFWNT9L_8tZ[249] , \b11_OFWNT9L_8tZ[248] , 
        \b11_OFWNT9L_8tZ[247] , \b11_OFWNT9L_8tZ[246] , 
        \b11_OFWNT9L_8tZ[245] , \b11_OFWNT9L_8tZ[244] , 
        \b11_OFWNT9L_8tZ[243] , \b11_OFWNT9L_8tZ[242] , 
        \b11_OFWNT9L_8tZ[241] , \b11_OFWNT9L_8tZ[240] , 
        \b11_OFWNT9L_8tZ[239] , \b11_OFWNT9L_8tZ[238] , 
        \b11_OFWNT9L_8tZ[237] , \b11_OFWNT9L_8tZ[236] , 
        \b11_OFWNT9L_8tZ[235] , \b11_OFWNT9L_8tZ[234] , 
        \b11_OFWNT9L_8tZ[233] , \b11_OFWNT9L_8tZ[232] , 
        \b11_OFWNT9L_8tZ[231] , \b11_OFWNT9L_8tZ[230] , 
        \b11_OFWNT9L_8tZ[229] , \b11_OFWNT9L_8tZ[228] , 
        \b11_OFWNT9L_8tZ[227] , \b11_OFWNT9L_8tZ[226] , 
        \b11_OFWNT9L_8tZ[225] , \b11_OFWNT9L_8tZ[224] , 
        \b11_OFWNT9L_8tZ[223] , \b11_OFWNT9L_8tZ[222] , 
        \b11_OFWNT9L_8tZ[221] , \b11_OFWNT9L_8tZ[220] , 
        \b11_OFWNT9L_8tZ[219] , \b11_OFWNT9L_8tZ[218] , 
        \b11_OFWNT9L_8tZ[217] , \b11_OFWNT9L_8tZ[216] , 
        \b11_OFWNT9L_8tZ[215] , \b11_OFWNT9L_8tZ[214] , 
        \b11_OFWNT9L_8tZ[213] , \b11_OFWNT9L_8tZ[212] , 
        \b11_OFWNT9L_8tZ[211] , \b11_OFWNT9L_8tZ[210] , 
        \b11_OFWNT9L_8tZ[209] , \b11_OFWNT9L_8tZ[208] , 
        \b11_OFWNT9L_8tZ[207] , \b11_OFWNT9L_8tZ[206] , 
        \b11_OFWNT9L_8tZ[205] , \b11_OFWNT9L_8tZ[204] , 
        \b11_OFWNT9L_8tZ[203] , \b11_OFWNT9L_8tZ[202] , 
        \b11_OFWNT9L_8tZ[201] , \b11_OFWNT9L_8tZ[200] , 
        \b11_OFWNT9L_8tZ[199] , \b11_OFWNT9L_8tZ[198] , 
        \b11_OFWNT9L_8tZ[197] , \b11_OFWNT9L_8tZ[196] , 
        \b11_OFWNT9L_8tZ[195] , \b11_OFWNT9L_8tZ[194] , 
        \b11_OFWNT9L_8tZ[193] , \b11_OFWNT9L_8tZ[192] , 
        \b11_OFWNT9L_8tZ[191] , \b11_OFWNT9L_8tZ[190] , 
        \b11_OFWNT9L_8tZ[189] , \b11_OFWNT9L_8tZ[188] , 
        \b11_OFWNT9L_8tZ[187] , \b11_OFWNT9L_8tZ[186] , 
        \b11_OFWNT9L_8tZ[185] , \b11_OFWNT9L_8tZ[184] , 
        \b11_OFWNT9L_8tZ[183] , \b11_OFWNT9L_8tZ[182] , 
        \b11_OFWNT9L_8tZ[181] , \b11_OFWNT9L_8tZ[180] , 
        \b11_OFWNT9L_8tZ[179] , \b11_OFWNT9L_8tZ[178] , 
        \b11_OFWNT9L_8tZ[177] , \b11_OFWNT9L_8tZ[176] , 
        \b11_OFWNT9L_8tZ[175] , \b11_OFWNT9L_8tZ[174] , 
        \b11_OFWNT9L_8tZ[173] , \b11_OFWNT9L_8tZ[172] , 
        \b11_OFWNT9L_8tZ[171] , \b11_OFWNT9L_8tZ[170] , 
        \b11_OFWNT9L_8tZ[169] , \b11_OFWNT9L_8tZ[168] , 
        \b11_OFWNT9L_8tZ[167] , \b11_OFWNT9L_8tZ[166] , 
        \b11_OFWNT9L_8tZ[165] , \b11_OFWNT9L_8tZ[164] , 
        \b11_OFWNT9L_8tZ[163] , \b11_OFWNT9L_8tZ[162] , 
        \b11_OFWNT9L_8tZ[161] , \b11_OFWNT9L_8tZ[160] , 
        \b11_OFWNT9L_8tZ[159] , \b11_OFWNT9L_8tZ[158] , 
        \b11_OFWNT9L_8tZ[157] , \b11_OFWNT9L_8tZ[156] , 
        \b11_OFWNT9L_8tZ[155] , \b11_OFWNT9L_8tZ[154] , 
        \b11_OFWNT9L_8tZ[153] , \b11_OFWNT9L_8tZ[152] , 
        \b11_OFWNT9L_8tZ[151] , \b11_OFWNT9L_8tZ[150] , 
        \b11_OFWNT9L_8tZ[149] , \b11_OFWNT9L_8tZ[148] , 
        \b11_OFWNT9L_8tZ[147] , \b11_OFWNT9L_8tZ[146] , 
        \b11_OFWNT9L_8tZ[145] , \b11_OFWNT9L_8tZ[144] , 
        \b11_OFWNT9L_8tZ[143] , \b11_OFWNT9L_8tZ[142] , 
        \b11_OFWNT9L_8tZ[141] , \b11_OFWNT9L_8tZ[140] , 
        \b11_OFWNT9L_8tZ[139] , \b11_OFWNT9L_8tZ[138] , 
        \b11_OFWNT9L_8tZ[137] , \b11_OFWNT9L_8tZ[136] , 
        \b11_OFWNT9L_8tZ[135] , \b11_OFWNT9L_8tZ[134] , 
        \b11_OFWNT9L_8tZ[133] , \b11_OFWNT9L_8tZ[132] , 
        \b11_OFWNT9L_8tZ[131] , \b11_OFWNT9L_8tZ[130] , 
        \b11_OFWNT9L_8tZ[129] , \b11_OFWNT9L_8tZ[128] , 
        \b11_OFWNT9L_8tZ[127] , \b11_OFWNT9L_8tZ[126] , 
        \b11_OFWNT9L_8tZ[125] , \b11_OFWNT9L_8tZ[124] , 
        \b11_OFWNT9L_8tZ[123] , \b11_OFWNT9L_8tZ[122] , 
        \b11_OFWNT9L_8tZ[121] , \b11_OFWNT9L_8tZ[120] , 
        \b11_OFWNT9L_8tZ[119] , \b11_OFWNT9L_8tZ[118] , 
        \b11_OFWNT9L_8tZ[117] , \b11_OFWNT9L_8tZ[116] , 
        \b11_OFWNT9L_8tZ[115] , \b11_OFWNT9L_8tZ[114] , 
        \b11_OFWNT9L_8tZ[113] , \b11_OFWNT9L_8tZ[112] , 
        \b11_OFWNT9L_8tZ[111] , \b11_OFWNT9L_8tZ[110] , 
        \b11_OFWNT9L_8tZ[109] , \b11_OFWNT9L_8tZ[108] , 
        \b11_OFWNT9L_8tZ[107] , \b11_OFWNT9L_8tZ[106] , 
        \b11_OFWNT9L_8tZ[105] , \b11_OFWNT9L_8tZ[104] , 
        \b11_OFWNT9L_8tZ[103] , \b11_OFWNT9L_8tZ[102] , 
        \b11_OFWNT9L_8tZ[101] , \b11_OFWNT9L_8tZ[100] , 
        \b11_OFWNT9L_8tZ[99] , \b11_OFWNT9L_8tZ[98] , 
        \b11_OFWNT9L_8tZ[97] , \b11_OFWNT9L_8tZ[96] , 
        \b11_OFWNT9L_8tZ[95] , \b11_OFWNT9L_8tZ[94] , 
        \b11_OFWNT9L_8tZ[93] , \b11_OFWNT9L_8tZ[92] , 
        \b11_OFWNT9L_8tZ[91] , \b11_OFWNT9L_8tZ[90] , 
        \b11_OFWNT9L_8tZ[89] , \b11_OFWNT9L_8tZ[88] , 
        \b11_OFWNT9L_8tZ[87] , \b11_OFWNT9L_8tZ[86] , 
        \b11_OFWNT9L_8tZ[85] , \b11_OFWNT9L_8tZ[84] , 
        \b11_OFWNT9L_8tZ[83] , \b11_OFWNT9L_8tZ[82] , 
        \b11_OFWNT9L_8tZ[81] , \b11_OFWNT9L_8tZ[80] , 
        \b11_OFWNT9L_8tZ[79] , \b11_OFWNT9L_8tZ[78] , 
        \b11_OFWNT9L_8tZ[77] , \b11_OFWNT9L_8tZ[76] , 
        \b11_OFWNT9L_8tZ[75] , \b11_OFWNT9L_8tZ[74] , 
        \b11_OFWNT9L_8tZ[73] , \b11_OFWNT9L_8tZ[72] , 
        \b11_OFWNT9L_8tZ[71] , \b11_OFWNT9L_8tZ[70] , 
        \b11_OFWNT9L_8tZ[69] , \b11_OFWNT9L_8tZ[68] , 
        \b11_OFWNT9L_8tZ[67] , \b11_OFWNT9L_8tZ[66] , 
        \b11_OFWNT9L_8tZ[65] , \b11_OFWNT9L_8tZ[64] , 
        \b11_OFWNT9L_8tZ[63] , \b11_OFWNT9L_8tZ[62] , 
        \b11_OFWNT9L_8tZ[61] , \b11_OFWNT9L_8tZ[60] , 
        \b11_OFWNT9L_8tZ[59] , \b11_OFWNT9L_8tZ[58] , 
        \b11_OFWNT9L_8tZ[57] , \b11_OFWNT9L_8tZ[56] , 
        \b11_OFWNT9L_8tZ[55] , \b11_OFWNT9L_8tZ[54] , 
        \b11_OFWNT9L_8tZ[53] , \b11_OFWNT9L_8tZ[52] , 
        \b11_OFWNT9L_8tZ[51] , \b11_OFWNT9L_8tZ[50] , 
        \b11_OFWNT9L_8tZ[49] , \b11_OFWNT9L_8tZ[48] , 
        \b11_OFWNT9L_8tZ[47] , \b11_OFWNT9L_8tZ[46] , 
        \b11_OFWNT9L_8tZ[45] , \b11_OFWNT9L_8tZ[44] , 
        \b11_OFWNT9L_8tZ[43] , \b11_OFWNT9L_8tZ[42] , 
        \b11_OFWNT9L_8tZ[41] , \b11_OFWNT9L_8tZ[40] , 
        \b11_OFWNT9L_8tZ[39] , \b11_OFWNT9L_8tZ[38] , 
        \b11_OFWNT9L_8tZ[37] , \b11_OFWNT9L_8tZ[36] , 
        \b11_OFWNT9L_8tZ[35] , \b11_OFWNT9L_8tZ[34] , 
        \b11_OFWNT9L_8tZ[33] , \b11_OFWNT9L_8tZ[32] , 
        \b11_OFWNT9L_8tZ[31] , \b11_OFWNT9L_8tZ[30] , 
        \b11_OFWNT9L_8tZ[29] , \b11_OFWNT9L_8tZ[28] , 
        \b11_OFWNT9L_8tZ[27] , \b11_OFWNT9L_8tZ[26] , 
        \b11_OFWNT9L_8tZ[25] , \b11_OFWNT9L_8tZ[24] , 
        \b11_OFWNT9L_8tZ[23] , \b11_OFWNT9L_8tZ[22] , 
        \b11_OFWNT9L_8tZ[21] , \b11_OFWNT9L_8tZ[20] , 
        \b11_OFWNT9L_8tZ[19] , \b11_OFWNT9L_8tZ[18] , 
        \b11_OFWNT9L_8tZ[17] , \b11_OFWNT9L_8tZ[16] , 
        \b11_OFWNT9L_8tZ[15] , \b11_OFWNT9L_8tZ[14] , 
        \b11_OFWNT9L_8tZ[13] , \b11_OFWNT9L_8tZ[12] , 
        \b11_OFWNT9L_8tZ[11] , \b11_OFWNT9L_8tZ[10] , 
        \b11_OFWNT9L_8tZ[9] , \b11_OFWNT9L_8tZ[8] , 
        \b11_OFWNT9L_8tZ[7] , \b11_OFWNT9L_8tZ[6] , 
        \b11_OFWNT9L_8tZ[5] , \b11_OFWNT9L_8tZ[4] , 
        \b11_OFWNT9L_8tZ[3] , \b11_OFWNT9L_8tZ[2] , 
        \b11_OFWNT9L_8tZ[1] , \b11_OFWNT9L_8tZ[0] }), .b8_SoWGfWYY(
        b8_SoWGfWYY), .b8_SoWGfWYY_i(b8_SoWGfWYY_i), .BW_clk_c(
        BW_clk_c), .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh), 
        .b11_PSyil9s_FMZ(b11_PSyil9s_FMZ), .b11_uRrc2XfY_XH(
        b11_uRrc2XfY_XH), .b4_PLyF(b4_PLyF), .b13_nUTQBgfDb_Z4D(
        b13_nUTQBgfDb_Z4D), .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), 
        .b16_nYhI39swMeEd_A78(b16_nYhI39swMeEd_A78), 
        .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), .b12_vABZ3qsY_Lyh(
        b12_vABZ3qsY_Lyh), .b11_vABZ3qsY_XH(b11_vABZ3qsY_XH), 
        .b7_PSyi3wy(b7_PSyi3wy), .b8_PSyiBgYG(b8_PSyiBgYG));
    SLE \mdiclink_reg[263]  (.D(temp1[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[263]_net_1 ));
    SLE \mdiclink_reg[344]  (.D(temp_so_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[344]_net_1 ));
    SLE \mdiclink_reg[307]  (.D(temp_count[30]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[307]_net_1 ));
    SLE \mdiclink_reg[289]  (.D(temp3[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[289]_net_1 ));
    SLE \mdiclink_reg[311]  (.D(temp_count[26]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[311]_net_1 ));
    SLE \mdiclink_reg[364]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[364]_net_1 ));
    SLE \mdiclink_reg[192]  (.D(fpga_shift_2[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[192]_net_1 ));
    SLE \mdiclink_reg[109]  (.D(\data_from_adc[4] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[109]_net_1 ));
    SLE \mdiclink_reg[239]  (.D(freq_6), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[239]_net_1 ));
    SLE \mdiclink_reg[181]  (.D(fpga_count[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[181]_net_1 ));
    SLE \mdiclink_reg[353]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[353]_net_1 ));
    SLE \mdiclink_reg[59]  (.D(\data_from_adc[8] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[59]_net_1 ));
    SLE \mdiclink_reg[178]  (.D(fpga_count[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[178]_net_1 ));
    SLE \mdiclink_reg[23]  (.D(BW_out_c[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[23]_net_1 ));
    SLE \mdiclink_reg[6]  (.D(BW_c[8]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[6]_net_1 ));
    SLE \mdiclink_reg[278]  (.D(temp2[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[278]_net_1 ));
    SLE \mdiclink_reg[124]  (.D(\data_from_adc[2] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[124]_net_1 ));
    SLE \mdiclink_reg[274]  (.D(temp2[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[274]_net_1 ));
    SLE \mdiclink_reg[11]  (.D(BW_c[3]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[11]_net_1 ));
    SLE \mdiclink_reg[325]  (.D(temp_count[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[325]_net_1 ));
    SLE \mdiclink_reg[143]  (.D(\data_from_adc[1] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[143]_net_1 ));
    SLE \mdiclink_reg[131]  (.D(\data_from_adc[2] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[131]_net_1 ));
    SLE \mdiclink_reg[312]  (.D(temp_count[25]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[312]_net_1 ));
    SLE \mdiclink_reg[9]  (.D(BW_c[5]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[9]_net_1 ));
    SLE \mdiclink_reg[273]  (.D(temp2[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[273]_net_1 ));
    SLE \mdiclink_reg[28]  (.D(BW_out_c[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[28]_net_1 ));
    SLE \mdiclink_reg[163]  (.D(dds_cos[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[163]_net_1 ));
    SLE \mdiclink_reg[107]  (.D(\data_from_adc[4] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[107]_net_1 ));
    SLE \mdiclink_reg[221]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[221]_net_1 ));
    SLE \mdiclink_reg[290]  (.D(temp3[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[290]_net_1 ));
    SLE \mdiclink_reg[106]  (.D(\data_from_adc[4] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[106]_net_1 ));
    SLE \mdiclink_reg[338]  (.D(temp_count_data[4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[338]_net_1 ));
    SLE \mdiclink_reg[100]  (.D(\data_from_adc[4] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[100]_net_1 ));
    SLE \mdiclink_reg[212]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[212]_net_1 ));
    SLE \mdiclink_reg[182]  (.D(fpga_count[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[182]_net_1 ));
    SLE \mdiclink_reg[26]  (.D(BW_out_c[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[26]_net_1 ));
    SLE \mdiclink_reg[374]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[374]_net_1 ));
    SLE \mdiclink_reg[71]  (.D(\data_from_adc[7] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[71]_net_1 ));
    SLE \mdiclink_reg[309]  (.D(temp_count[28]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[309]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \mdiclink_reg[321]  (.D(temp_count[16]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[321]_net_1 ));
    SLE \mdiclink_reg[206]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[206]_net_1 ));
    SLE \mdiclink_reg[55]  (.D(\data_from_adc[8] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[55]_net_1 ));
    SLE \mdiclink_reg[217]  (.D(fr_adc_count[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[217]_net_1 ));
    SLE \mdiclink_reg[13]  (.D(BW_c[1]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[13]_net_1 ));
    SLE \mdiclink_reg[132]  (.D(\data_from_adc[2] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[132]_net_1 ));
    SLE \mdiclink_reg[62]  (.D(\data_from_adc[7] [11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[62]_net_1 ));
    SLE \mdiclink_reg[145]  (.D(\data_from_adc[1] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[145]_net_1 ));
    SLE \mdiclink_reg[154]  (.D(\data_from_adc[0] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[154]_net_1 ));
    SLE \mdiclink_reg[300]  (.D(temp3[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[300]_net_1 ));
    SLE \mdiclink_reg[355]  (.D(freq_14), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[355]_net_1 ));
    SLE \mdiclink_reg[165]  (.D(dds_cos[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[165]_net_1 ));
    SLE \mdiclink_reg[336]  (.D(temp_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[336]_net_1 ));
    SLE \mdiclink_reg[295]  (.D(temp3[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[295]_net_1 ));
    SLE \mdiclink_reg[280]  (.D(temp2[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[280]_net_1 ));
    SLE \mdiclink_reg[18]  (.D(BW_out_c[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[18]_net_1 ));
    SLE \mdiclink_reg[173]  (.D(dds_sin[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[173]_net_1 ));
    SLE \mdiclink_reg[8]  (.D(BW_c[6]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[8]_net_1 ));
    SLE \mdiclink_reg[50]  (.D(\data_from_adc[8] [11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[50]_net_1 ));
    SLE \mdiclink_reg[251]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[251]_net_1 ));
    SLE \mdiclink_reg[73]  (.D(\data_from_adc[7] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[73]_net_1 ));
    SLE \mdiclink_reg[322]  (.D(temp_count[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[322]_net_1 ));
    SLE \mdiclink_reg[16]  (.D(BW_out_c[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[16]_net_1 ));
    SLE \mdiclink_reg[64]  (.D(\data_from_adc[7] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[64]_net_1 ));
    SLE \mdiclink_reg[57]  (.D(\data_from_adc[8] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[57]_net_1 ));
    SLE \mdiclink_reg[230]  (.D(freq_15), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[230]_net_1 ));
    SLE \mdiclink_reg[351]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[351]_net_1 ));
    SLE \mdiclink_reg[222]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[222]_net_1 ));
    SLE \mdiclink_reg[347]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[347]_net_1 ));
    SLE \mdiclink_reg[78]  (.D(\data_from_adc[6] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[78]_net_1 ));
    SLE \mdiclink_reg[285]  (.D(temp2[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[285]_net_1 ));
    SLE \mdiclink_reg[367]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[367]_net_1 ));
    SLE \mdiclink_reg[303]  (.D(temp3[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[303]_net_1 ));
    SLE \mdiclink_reg[227]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[227]_net_1 ));
    SLE \mdiclink_reg[32]  (.D(dac1_db_c[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[32]_net_1 ));
    SLE \mdiclink_reg[149]  (.D(\data_from_adc[0] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[149]_net_1 ));
    SLE \mdiclink_reg[76]  (.D(\data_from_adc[6] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[76]_net_1 ));
    SLE \mdiclink_reg[175]  (.D(fpga_count[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[175]_net_1 ));
    SLE \mdiclink_reg[219]  (.D(fr_adc_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[219]_net_1 ));
    SLE \mdiclink_reg[235]  (.D(freq_10), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[235]_net_1 ));
    SLE \mdiclink_reg[169]  (.D(dds_sin[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[169]_net_1 ));
    b11_OFWNT9s_8tZ_Z2_x b3_SoW_0 (.b11_OFWNT9L_8tZ({
        \b11_OFWNT9L_8tZ[376] , \b11_OFWNT9L_8tZ[375] , 
        \b11_OFWNT9L_8tZ[374] , \b11_OFWNT9L_8tZ[373] , 
        \b11_OFWNT9L_8tZ[372] , \b11_OFWNT9L_8tZ[371] , 
        \b11_OFWNT9L_8tZ[370] , \b11_OFWNT9L_8tZ[369] , 
        \b11_OFWNT9L_8tZ[368] , \b11_OFWNT9L_8tZ[367] , 
        \b11_OFWNT9L_8tZ[366] , \b11_OFWNT9L_8tZ[365] , 
        \b11_OFWNT9L_8tZ[364] , \b11_OFWNT9L_8tZ[363] , 
        \b11_OFWNT9L_8tZ[362] , \b11_OFWNT9L_8tZ[361] , 
        \b11_OFWNT9L_8tZ[360] , \b11_OFWNT9L_8tZ[359] , 
        \b11_OFWNT9L_8tZ[358] , \b11_OFWNT9L_8tZ[357] , 
        \b11_OFWNT9L_8tZ[356] , \b11_OFWNT9L_8tZ[355] , 
        \b11_OFWNT9L_8tZ[354] , \b11_OFWNT9L_8tZ[353] , 
        \b11_OFWNT9L_8tZ[352] , \b11_OFWNT9L_8tZ[351] , 
        \b11_OFWNT9L_8tZ[350] , \b11_OFWNT9L_8tZ[349] , 
        \b11_OFWNT9L_8tZ[348] , \b11_OFWNT9L_8tZ[347] , 
        \b11_OFWNT9L_8tZ[346] , \b11_OFWNT9L_8tZ[345] , 
        \b11_OFWNT9L_8tZ[344] , \b11_OFWNT9L_8tZ[343] , 
        \b11_OFWNT9L_8tZ[342] , \b11_OFWNT9L_8tZ[341] , 
        \b11_OFWNT9L_8tZ[340] , \b11_OFWNT9L_8tZ[339] , 
        \b11_OFWNT9L_8tZ[338] , \b11_OFWNT9L_8tZ[337] , 
        \b11_OFWNT9L_8tZ[336] , \b11_OFWNT9L_8tZ[335] , 
        \b11_OFWNT9L_8tZ[334] , \b11_OFWNT9L_8tZ[333] , 
        \b11_OFWNT9L_8tZ[332] , \b11_OFWNT9L_8tZ[331] , 
        \b11_OFWNT9L_8tZ[330] , \b11_OFWNT9L_8tZ[329] , 
        \b11_OFWNT9L_8tZ[328] , \b11_OFWNT9L_8tZ[327] , 
        \b11_OFWNT9L_8tZ[326] , \b11_OFWNT9L_8tZ[325] , 
        \b11_OFWNT9L_8tZ[324] , \b11_OFWNT9L_8tZ[323] , 
        \b11_OFWNT9L_8tZ[322] , \b11_OFWNT9L_8tZ[321] , 
        \b11_OFWNT9L_8tZ[320] , \b11_OFWNT9L_8tZ[319] , 
        \b11_OFWNT9L_8tZ[318] , \b11_OFWNT9L_8tZ[317] , 
        \b11_OFWNT9L_8tZ[316] , \b11_OFWNT9L_8tZ[315] , 
        \b11_OFWNT9L_8tZ[314] , \b11_OFWNT9L_8tZ[313] , 
        \b11_OFWNT9L_8tZ[312] , \b11_OFWNT9L_8tZ[311] , 
        \b11_OFWNT9L_8tZ[310] , \b11_OFWNT9L_8tZ[309] , 
        \b11_OFWNT9L_8tZ[308] , \b11_OFWNT9L_8tZ[307] , 
        \b11_OFWNT9L_8tZ[306] , \b11_OFWNT9L_8tZ[305] , 
        \b11_OFWNT9L_8tZ[304] , \b11_OFWNT9L_8tZ[303] , 
        \b11_OFWNT9L_8tZ[302] , \b11_OFWNT9L_8tZ[301] , 
        \b11_OFWNT9L_8tZ[300] , \b11_OFWNT9L_8tZ[299] , 
        \b11_OFWNT9L_8tZ[298] , \b11_OFWNT9L_8tZ[297] , 
        \b11_OFWNT9L_8tZ[296] , \b11_OFWNT9L_8tZ[295] , 
        \b11_OFWNT9L_8tZ[294] , \b11_OFWNT9L_8tZ[293] , 
        \b11_OFWNT9L_8tZ[292] , \b11_OFWNT9L_8tZ[291] , 
        \b11_OFWNT9L_8tZ[290] , \b11_OFWNT9L_8tZ[289] , 
        \b11_OFWNT9L_8tZ[288] , \b11_OFWNT9L_8tZ[287] , 
        \b11_OFWNT9L_8tZ[286] , \b11_OFWNT9L_8tZ[285] , 
        \b11_OFWNT9L_8tZ[284] , \b11_OFWNT9L_8tZ[283] , 
        \b11_OFWNT9L_8tZ[282] , \b11_OFWNT9L_8tZ[281] , 
        \b11_OFWNT9L_8tZ[280] , \b11_OFWNT9L_8tZ[279] , 
        \b11_OFWNT9L_8tZ[278] , \b11_OFWNT9L_8tZ[277] , 
        \b11_OFWNT9L_8tZ[276] , \b11_OFWNT9L_8tZ[275] , 
        \b11_OFWNT9L_8tZ[274] , \b11_OFWNT9L_8tZ[273] , 
        \b11_OFWNT9L_8tZ[272] , \b11_OFWNT9L_8tZ[271] , 
        \b11_OFWNT9L_8tZ[270] , \b11_OFWNT9L_8tZ[269] , 
        \b11_OFWNT9L_8tZ[268] , \b11_OFWNT9L_8tZ[267] , 
        \b11_OFWNT9L_8tZ[266] , \b11_OFWNT9L_8tZ[265] , 
        \b11_OFWNT9L_8tZ[264] , \b11_OFWNT9L_8tZ[263] , 
        \b11_OFWNT9L_8tZ[262] , \b11_OFWNT9L_8tZ[261] , 
        \b11_OFWNT9L_8tZ[260] , \b11_OFWNT9L_8tZ[259] , 
        \b11_OFWNT9L_8tZ[258] , \b11_OFWNT9L_8tZ[257] , 
        \b11_OFWNT9L_8tZ[256] , \b11_OFWNT9L_8tZ[255] , 
        \b11_OFWNT9L_8tZ[254] , \b11_OFWNT9L_8tZ[253] , 
        \b11_OFWNT9L_8tZ[252] , \b11_OFWNT9L_8tZ[251] , 
        \b11_OFWNT9L_8tZ[250] , \b11_OFWNT9L_8tZ[249] , 
        \b11_OFWNT9L_8tZ[248] , \b11_OFWNT9L_8tZ[247] , 
        \b11_OFWNT9L_8tZ[246] , \b11_OFWNT9L_8tZ[245] , 
        \b11_OFWNT9L_8tZ[244] , \b11_OFWNT9L_8tZ[243] , 
        \b11_OFWNT9L_8tZ[242] , \b11_OFWNT9L_8tZ[241] , 
        \b11_OFWNT9L_8tZ[240] , \b11_OFWNT9L_8tZ[239] , 
        \b11_OFWNT9L_8tZ[238] , \b11_OFWNT9L_8tZ[237] , 
        \b11_OFWNT9L_8tZ[236] , \b11_OFWNT9L_8tZ[235] , 
        \b11_OFWNT9L_8tZ[234] , \b11_OFWNT9L_8tZ[233] , 
        \b11_OFWNT9L_8tZ[232] , \b11_OFWNT9L_8tZ[231] , 
        \b11_OFWNT9L_8tZ[230] , \b11_OFWNT9L_8tZ[229] , 
        \b11_OFWNT9L_8tZ[228] , \b11_OFWNT9L_8tZ[227] , 
        \b11_OFWNT9L_8tZ[226] , \b11_OFWNT9L_8tZ[225] , 
        \b11_OFWNT9L_8tZ[224] , \b11_OFWNT9L_8tZ[223] , 
        \b11_OFWNT9L_8tZ[222] , \b11_OFWNT9L_8tZ[221] , 
        \b11_OFWNT9L_8tZ[220] , \b11_OFWNT9L_8tZ[219] , 
        \b11_OFWNT9L_8tZ[218] , \b11_OFWNT9L_8tZ[217] , 
        \b11_OFWNT9L_8tZ[216] , \b11_OFWNT9L_8tZ[215] , 
        \b11_OFWNT9L_8tZ[214] , \b11_OFWNT9L_8tZ[213] , 
        \b11_OFWNT9L_8tZ[212] , \b11_OFWNT9L_8tZ[211] , 
        \b11_OFWNT9L_8tZ[210] , \b11_OFWNT9L_8tZ[209] , 
        \b11_OFWNT9L_8tZ[208] , \b11_OFWNT9L_8tZ[207] , 
        \b11_OFWNT9L_8tZ[206] , \b11_OFWNT9L_8tZ[205] , 
        \b11_OFWNT9L_8tZ[204] , \b11_OFWNT9L_8tZ[203] , 
        \b11_OFWNT9L_8tZ[202] , \b11_OFWNT9L_8tZ[201] , 
        \b11_OFWNT9L_8tZ[200] , \b11_OFWNT9L_8tZ[199] , 
        \b11_OFWNT9L_8tZ[198] , \b11_OFWNT9L_8tZ[197] , 
        \b11_OFWNT9L_8tZ[196] , \b11_OFWNT9L_8tZ[195] , 
        \b11_OFWNT9L_8tZ[194] , \b11_OFWNT9L_8tZ[193] , 
        \b11_OFWNT9L_8tZ[192] , \b11_OFWNT9L_8tZ[191] , 
        \b11_OFWNT9L_8tZ[190] , \b11_OFWNT9L_8tZ[189] , 
        \b11_OFWNT9L_8tZ[188] , \b11_OFWNT9L_8tZ[187] , 
        \b11_OFWNT9L_8tZ[186] , \b11_OFWNT9L_8tZ[185] , 
        \b11_OFWNT9L_8tZ[184] , \b11_OFWNT9L_8tZ[183] , 
        \b11_OFWNT9L_8tZ[182] , \b11_OFWNT9L_8tZ[181] , 
        \b11_OFWNT9L_8tZ[180] , \b11_OFWNT9L_8tZ[179] , 
        \b11_OFWNT9L_8tZ[178] , \b11_OFWNT9L_8tZ[177] , 
        \b11_OFWNT9L_8tZ[176] , \b11_OFWNT9L_8tZ[175] , 
        \b11_OFWNT9L_8tZ[174] , \b11_OFWNT9L_8tZ[173] , 
        \b11_OFWNT9L_8tZ[172] , \b11_OFWNT9L_8tZ[171] , 
        \b11_OFWNT9L_8tZ[170] , \b11_OFWNT9L_8tZ[169] , 
        \b11_OFWNT9L_8tZ[168] , \b11_OFWNT9L_8tZ[167] , 
        \b11_OFWNT9L_8tZ[166] , \b11_OFWNT9L_8tZ[165] , 
        \b11_OFWNT9L_8tZ[164] , \b11_OFWNT9L_8tZ[163] , 
        \b11_OFWNT9L_8tZ[162] , \b11_OFWNT9L_8tZ[161] , 
        \b11_OFWNT9L_8tZ[160] , \b11_OFWNT9L_8tZ[159] , 
        \b11_OFWNT9L_8tZ[158] , \b11_OFWNT9L_8tZ[157] , 
        \b11_OFWNT9L_8tZ[156] , \b11_OFWNT9L_8tZ[155] , 
        \b11_OFWNT9L_8tZ[154] , \b11_OFWNT9L_8tZ[153] , 
        \b11_OFWNT9L_8tZ[152] , \b11_OFWNT9L_8tZ[151] , 
        \b11_OFWNT9L_8tZ[150] , \b11_OFWNT9L_8tZ[149] , 
        \b11_OFWNT9L_8tZ[148] , \b11_OFWNT9L_8tZ[147] , 
        \b11_OFWNT9L_8tZ[146] , \b11_OFWNT9L_8tZ[145] , 
        \b11_OFWNT9L_8tZ[144] , \b11_OFWNT9L_8tZ[143] , 
        \b11_OFWNT9L_8tZ[142] , \b11_OFWNT9L_8tZ[141] , 
        \b11_OFWNT9L_8tZ[140] , \b11_OFWNT9L_8tZ[139] , 
        \b11_OFWNT9L_8tZ[138] , \b11_OFWNT9L_8tZ[137] , 
        \b11_OFWNT9L_8tZ[136] , \b11_OFWNT9L_8tZ[135] , 
        \b11_OFWNT9L_8tZ[134] , \b11_OFWNT9L_8tZ[133] , 
        \b11_OFWNT9L_8tZ[132] , \b11_OFWNT9L_8tZ[131] , 
        \b11_OFWNT9L_8tZ[130] , \b11_OFWNT9L_8tZ[129] , 
        \b11_OFWNT9L_8tZ[128] , \b11_OFWNT9L_8tZ[127] , 
        \b11_OFWNT9L_8tZ[126] , \b11_OFWNT9L_8tZ[125] , 
        \b11_OFWNT9L_8tZ[124] , \b11_OFWNT9L_8tZ[123] , 
        \b11_OFWNT9L_8tZ[122] , \b11_OFWNT9L_8tZ[121] , 
        \b11_OFWNT9L_8tZ[120] , \b11_OFWNT9L_8tZ[119] , 
        \b11_OFWNT9L_8tZ[118] , \b11_OFWNT9L_8tZ[117] , 
        \b11_OFWNT9L_8tZ[116] , \b11_OFWNT9L_8tZ[115] , 
        \b11_OFWNT9L_8tZ[114] , \b11_OFWNT9L_8tZ[113] , 
        \b11_OFWNT9L_8tZ[112] , \b11_OFWNT9L_8tZ[111] , 
        \b11_OFWNT9L_8tZ[110] , \b11_OFWNT9L_8tZ[109] , 
        \b11_OFWNT9L_8tZ[108] , \b11_OFWNT9L_8tZ[107] , 
        \b11_OFWNT9L_8tZ[106] , \b11_OFWNT9L_8tZ[105] , 
        \b11_OFWNT9L_8tZ[104] , \b11_OFWNT9L_8tZ[103] , 
        \b11_OFWNT9L_8tZ[102] , \b11_OFWNT9L_8tZ[101] , 
        \b11_OFWNT9L_8tZ[100] , \b11_OFWNT9L_8tZ[99] , 
        \b11_OFWNT9L_8tZ[98] , \b11_OFWNT9L_8tZ[97] , 
        \b11_OFWNT9L_8tZ[96] , \b11_OFWNT9L_8tZ[95] , 
        \b11_OFWNT9L_8tZ[94] , \b11_OFWNT9L_8tZ[93] , 
        \b11_OFWNT9L_8tZ[92] , \b11_OFWNT9L_8tZ[91] , 
        \b11_OFWNT9L_8tZ[90] , \b11_OFWNT9L_8tZ[89] , 
        \b11_OFWNT9L_8tZ[88] , \b11_OFWNT9L_8tZ[87] , 
        \b11_OFWNT9L_8tZ[86] , \b11_OFWNT9L_8tZ[85] , 
        \b11_OFWNT9L_8tZ[84] , \b11_OFWNT9L_8tZ[83] , 
        \b11_OFWNT9L_8tZ[82] , \b11_OFWNT9L_8tZ[81] , 
        \b11_OFWNT9L_8tZ[80] , \b11_OFWNT9L_8tZ[79] , 
        \b11_OFWNT9L_8tZ[78] , \b11_OFWNT9L_8tZ[77] , 
        \b11_OFWNT9L_8tZ[76] , \b11_OFWNT9L_8tZ[75] , 
        \b11_OFWNT9L_8tZ[74] , \b11_OFWNT9L_8tZ[73] , 
        \b11_OFWNT9L_8tZ[72] , \b11_OFWNT9L_8tZ[71] , 
        \b11_OFWNT9L_8tZ[70] , \b11_OFWNT9L_8tZ[69] , 
        \b11_OFWNT9L_8tZ[68] , \b11_OFWNT9L_8tZ[67] , 
        \b11_OFWNT9L_8tZ[66] , \b11_OFWNT9L_8tZ[65] , 
        \b11_OFWNT9L_8tZ[64] , \b11_OFWNT9L_8tZ[63] , 
        \b11_OFWNT9L_8tZ[62] , \b11_OFWNT9L_8tZ[61] , 
        \b11_OFWNT9L_8tZ[60] , \b11_OFWNT9L_8tZ[59] , 
        \b11_OFWNT9L_8tZ[58] , \b11_OFWNT9L_8tZ[57] , 
        \b11_OFWNT9L_8tZ[56] , \b11_OFWNT9L_8tZ[55] , 
        \b11_OFWNT9L_8tZ[54] , \b11_OFWNT9L_8tZ[53] , 
        \b11_OFWNT9L_8tZ[52] , \b11_OFWNT9L_8tZ[51] , 
        \b11_OFWNT9L_8tZ[50] , \b11_OFWNT9L_8tZ[49] , 
        \b11_OFWNT9L_8tZ[48] , \b11_OFWNT9L_8tZ[47] , 
        \b11_OFWNT9L_8tZ[46] , \b11_OFWNT9L_8tZ[45] , 
        \b11_OFWNT9L_8tZ[44] , \b11_OFWNT9L_8tZ[43] , 
        \b11_OFWNT9L_8tZ[42] , \b11_OFWNT9L_8tZ[41] , 
        \b11_OFWNT9L_8tZ[40] , \b11_OFWNT9L_8tZ[39] , 
        \b11_OFWNT9L_8tZ[38] , \b11_OFWNT9L_8tZ[37] , 
        \b11_OFWNT9L_8tZ[36] , \b11_OFWNT9L_8tZ[35] , 
        \b11_OFWNT9L_8tZ[34] , \b11_OFWNT9L_8tZ[33] , 
        \b11_OFWNT9L_8tZ[32] , \b11_OFWNT9L_8tZ[31] , 
        \b11_OFWNT9L_8tZ[30] , \b11_OFWNT9L_8tZ[29] , 
        \b11_OFWNT9L_8tZ[28] , \b11_OFWNT9L_8tZ[27] , 
        \b11_OFWNT9L_8tZ[26] , \b11_OFWNT9L_8tZ[25] , 
        \b11_OFWNT9L_8tZ[24] , \b11_OFWNT9L_8tZ[23] , 
        \b11_OFWNT9L_8tZ[22] , \b11_OFWNT9L_8tZ[21] , 
        \b11_OFWNT9L_8tZ[20] , \b11_OFWNT9L_8tZ[19] , 
        \b11_OFWNT9L_8tZ[18] , \b11_OFWNT9L_8tZ[17] , 
        \b11_OFWNT9L_8tZ[16] , \b11_OFWNT9L_8tZ[15] , 
        \b11_OFWNT9L_8tZ[14] , \b11_OFWNT9L_8tZ[13] , 
        \b11_OFWNT9L_8tZ[12] , \b11_OFWNT9L_8tZ[11] , 
        \b11_OFWNT9L_8tZ[10] , \b11_OFWNT9L_8tZ[9] , 
        \b11_OFWNT9L_8tZ[8] , \b11_OFWNT9L_8tZ[7] , 
        \b11_OFWNT9L_8tZ[6] , \b11_OFWNT9L_8tZ[5] , 
        \b11_OFWNT9L_8tZ[4] , \b11_OFWNT9L_8tZ[3] , 
        \b11_OFWNT9L_8tZ[2] , \b11_OFWNT9L_8tZ[1] , 
        \b11_OFWNT9L_8tZ[0] }), .mdiclink_reg({
        \mdiclink_reg[376]_net_1 , \mdiclink_reg[375]_net_1 , 
        \mdiclink_reg[374]_net_1 , \mdiclink_reg[373]_net_1 , 
        \mdiclink_reg[372]_net_1 , \mdiclink_reg[371]_net_1 , 
        \mdiclink_reg[370]_net_1 , \mdiclink_reg[369]_net_1 , 
        \mdiclink_reg[368]_net_1 , \mdiclink_reg[367]_net_1 , 
        \mdiclink_reg[366]_net_1 , \mdiclink_reg[365]_net_1 , 
        \mdiclink_reg[364]_net_1 , \mdiclink_reg[363]_net_1 , 
        \mdiclink_reg[362]_net_1 , \mdiclink_reg[361]_net_1 , 
        \mdiclink_reg[360]_net_1 , \mdiclink_reg[359]_net_1 , 
        \mdiclink_reg[358]_net_1 , \mdiclink_reg[357]_net_1 , 
        \mdiclink_reg[356]_net_1 , \mdiclink_reg[355]_net_1 , 
        \mdiclink_reg[354]_net_1 , \mdiclink_reg[353]_net_1 , 
        \mdiclink_reg[352]_net_1 , \mdiclink_reg[351]_net_1 , 
        \mdiclink_reg[350]_net_1 , \mdiclink_reg[349]_net_1 , 
        \mdiclink_reg[348]_net_1 , \mdiclink_reg[347]_net_1 , 
        \mdiclink_reg[346]_net_1 , \mdiclink_reg[345]_net_1 , 
        \mdiclink_reg[344]_net_1 , \mdiclink_reg[343]_net_1 , 
        \mdiclink_reg[342]_net_1 , \mdiclink_reg[341]_net_1 , 
        \mdiclink_reg[340]_net_1 , \mdiclink_reg[339]_net_1 , 
        \mdiclink_reg[338]_net_1 , \mdiclink_reg[337]_net_1 , 
        \mdiclink_reg[336]_net_1 , \mdiclink_reg[335]_net_1 , 
        \mdiclink_reg[334]_net_1 , \mdiclink_reg[333]_net_1 , 
        \mdiclink_reg[332]_net_1 , \mdiclink_reg[331]_net_1 , 
        \mdiclink_reg[330]_net_1 , \mdiclink_reg[329]_net_1 , 
        \mdiclink_reg[328]_net_1 , \mdiclink_reg[327]_net_1 , 
        \mdiclink_reg[326]_net_1 , \mdiclink_reg[325]_net_1 , 
        \mdiclink_reg[324]_net_1 , \mdiclink_reg[323]_net_1 , 
        \mdiclink_reg[322]_net_1 , \mdiclink_reg[321]_net_1 , 
        \mdiclink_reg[320]_net_1 , \mdiclink_reg[319]_net_1 , 
        \mdiclink_reg[318]_net_1 , \mdiclink_reg[317]_net_1 , 
        \mdiclink_reg[316]_net_1 , \mdiclink_reg[315]_net_1 , 
        \mdiclink_reg[314]_net_1 , \mdiclink_reg[313]_net_1 , 
        \mdiclink_reg[312]_net_1 , \mdiclink_reg[311]_net_1 , 
        \mdiclink_reg[310]_net_1 , \mdiclink_reg[309]_net_1 , 
        \mdiclink_reg[308]_net_1 , \mdiclink_reg[307]_net_1 , 
        \mdiclink_reg[306]_net_1 , \mdiclink_reg[305]_net_1 , 
        \mdiclink_reg[304]_net_1 , \mdiclink_reg[303]_net_1 , 
        \mdiclink_reg[302]_net_1 , \mdiclink_reg[301]_net_1 , 
        \mdiclink_reg[300]_net_1 , \mdiclink_reg[299]_net_1 , 
        \mdiclink_reg[298]_net_1 , \mdiclink_reg[297]_net_1 , 
        \mdiclink_reg[296]_net_1 , \mdiclink_reg[295]_net_1 , 
        \mdiclink_reg[294]_net_1 , \mdiclink_reg[293]_net_1 , 
        \mdiclink_reg[292]_net_1 , \mdiclink_reg[291]_net_1 , 
        \mdiclink_reg[290]_net_1 , \mdiclink_reg[289]_net_1 , 
        \mdiclink_reg[288]_net_1 , \mdiclink_reg[287]_net_1 , 
        \mdiclink_reg[286]_net_1 , \mdiclink_reg[285]_net_1 , 
        \mdiclink_reg[284]_net_1 , \mdiclink_reg[283]_net_1 , 
        \mdiclink_reg[282]_net_1 , \mdiclink_reg[281]_net_1 , 
        \mdiclink_reg[280]_net_1 , \mdiclink_reg[279]_net_1 , 
        \mdiclink_reg[278]_net_1 , \mdiclink_reg[277]_net_1 , 
        \mdiclink_reg[276]_net_1 , \mdiclink_reg[275]_net_1 , 
        \mdiclink_reg[274]_net_1 , \mdiclink_reg[273]_net_1 , 
        \mdiclink_reg[272]_net_1 , \mdiclink_reg[271]_net_1 , 
        \mdiclink_reg[270]_net_1 , \mdiclink_reg[269]_net_1 , 
        \mdiclink_reg[268]_net_1 , \mdiclink_reg[267]_net_1 , 
        \mdiclink_reg[266]_net_1 , \mdiclink_reg[265]_net_1 , 
        \mdiclink_reg[264]_net_1 , \mdiclink_reg[263]_net_1 , 
        \mdiclink_reg[262]_net_1 , \mdiclink_reg[261]_net_1 , 
        \mdiclink_reg[260]_net_1 , \mdiclink_reg[259]_net_1 , 
        \mdiclink_reg[258]_net_1 , \mdiclink_reg[257]_net_1 , 
        \mdiclink_reg[256]_net_1 , \mdiclink_reg[255]_net_1 , 
        \mdiclink_reg[254]_net_1 , \mdiclink_reg[253]_net_1 , 
        \mdiclink_reg[252]_net_1 , \mdiclink_reg[251]_net_1 , 
        \mdiclink_reg[250]_net_1 , \mdiclink_reg[249]_net_1 , 
        \mdiclink_reg[248]_net_1 , \mdiclink_reg[247]_net_1 , 
        \mdiclink_reg[246]_net_1 , \mdiclink_reg[245]_net_1 , 
        \mdiclink_reg[244]_net_1 , \mdiclink_reg[243]_net_1 , 
        \mdiclink_reg[242]_net_1 , \mdiclink_reg[241]_net_1 , 
        \mdiclink_reg[240]_net_1 , \mdiclink_reg[239]_net_1 , 
        \mdiclink_reg[238]_net_1 , \mdiclink_reg[237]_net_1 , 
        \mdiclink_reg[236]_net_1 , \mdiclink_reg[235]_net_1 , 
        \mdiclink_reg[234]_net_1 , \mdiclink_reg[233]_net_1 , 
        \mdiclink_reg[232]_net_1 , \mdiclink_reg[231]_net_1 , 
        \mdiclink_reg[230]_net_1 , \mdiclink_reg[229]_net_1 , 
        \mdiclink_reg[228]_net_1 , \mdiclink_reg[227]_net_1 , 
        \mdiclink_reg[226]_net_1 , \mdiclink_reg[225]_net_1 , 
        \mdiclink_reg[224]_net_1 , \mdiclink_reg[223]_net_1 , 
        \mdiclink_reg[222]_net_1 , \mdiclink_reg[221]_net_1 , 
        \mdiclink_reg[220]_net_1 , \mdiclink_reg[219]_net_1 , 
        \mdiclink_reg[218]_net_1 , \mdiclink_reg[217]_net_1 , 
        \mdiclink_reg[216]_net_1 , \mdiclink_reg[215]_net_1 , 
        \mdiclink_reg[214]_net_1 , \mdiclink_reg[213]_net_1 , 
        \mdiclink_reg[212]_net_1 , \mdiclink_reg[211]_net_1 , 
        \mdiclink_reg[210]_net_1 , \mdiclink_reg[209]_net_1 , 
        \mdiclink_reg[208]_net_1 , \mdiclink_reg[207]_net_1 , 
        \mdiclink_reg[206]_net_1 , \mdiclink_reg[205]_net_1 , 
        \mdiclink_reg[204]_net_1 , \mdiclink_reg[203]_net_1 , 
        \mdiclink_reg[202]_net_1 , \mdiclink_reg[201]_net_1 , 
        \mdiclink_reg[200]_net_1 , \mdiclink_reg[199]_net_1 , 
        \mdiclink_reg[198]_net_1 , \mdiclink_reg[197]_net_1 , 
        \mdiclink_reg[196]_net_1 , \mdiclink_reg[195]_net_1 , 
        \mdiclink_reg[194]_net_1 , \mdiclink_reg[193]_net_1 , 
        \mdiclink_reg[192]_net_1 , \mdiclink_reg[191]_net_1 , 
        \mdiclink_reg[190]_net_1 , \mdiclink_reg[189]_net_1 , 
        \mdiclink_reg[188]_net_1 , \mdiclink_reg[187]_net_1 , 
        \mdiclink_reg[186]_net_1 , \mdiclink_reg[185]_net_1 , 
        \mdiclink_reg[184]_net_1 , \mdiclink_reg[183]_net_1 , 
        \mdiclink_reg[182]_net_1 , \mdiclink_reg[181]_net_1 , 
        \mdiclink_reg[180]_net_1 , \mdiclink_reg[179]_net_1 , 
        \mdiclink_reg[178]_net_1 , \mdiclink_reg[177]_net_1 , 
        \mdiclink_reg[176]_net_1 , \mdiclink_reg[175]_net_1 , 
        \mdiclink_reg[174]_net_1 , \mdiclink_reg[173]_net_1 , 
        \mdiclink_reg[172]_net_1 , \mdiclink_reg[171]_net_1 , 
        \mdiclink_reg[170]_net_1 , \mdiclink_reg[169]_net_1 , 
        \mdiclink_reg[168]_net_1 , \mdiclink_reg[167]_net_1 , 
        \mdiclink_reg[166]_net_1 , \mdiclink_reg[165]_net_1 , 
        \mdiclink_reg[164]_net_1 , \mdiclink_reg[163]_net_1 , 
        \mdiclink_reg[162]_net_1 , \mdiclink_reg[161]_net_1 , 
        \mdiclink_reg[160]_net_1 , \mdiclink_reg[159]_net_1 , 
        \mdiclink_reg[158]_net_1 , \mdiclink_reg[157]_net_1 , 
        \mdiclink_reg[156]_net_1 , \mdiclink_reg[155]_net_1 , 
        \mdiclink_reg[154]_net_1 , \mdiclink_reg[153]_net_1 , 
        \mdiclink_reg[152]_net_1 , \mdiclink_reg[151]_net_1 , 
        \mdiclink_reg[150]_net_1 , \mdiclink_reg[149]_net_1 , 
        \mdiclink_reg[148]_net_1 , \mdiclink_reg[147]_net_1 , 
        \mdiclink_reg[146]_net_1 , \mdiclink_reg[145]_net_1 , 
        \mdiclink_reg[144]_net_1 , \mdiclink_reg[143]_net_1 , 
        \mdiclink_reg[142]_net_1 , \mdiclink_reg[141]_net_1 , 
        \mdiclink_reg[140]_net_1 , \mdiclink_reg[139]_net_1 , 
        \mdiclink_reg[138]_net_1 , \mdiclink_reg[137]_net_1 , 
        \mdiclink_reg[136]_net_1 , \mdiclink_reg[135]_net_1 , 
        \mdiclink_reg[134]_net_1 , \mdiclink_reg[133]_net_1 , 
        \mdiclink_reg[132]_net_1 , \mdiclink_reg[131]_net_1 , 
        \mdiclink_reg[130]_net_1 , \mdiclink_reg[129]_net_1 , 
        \mdiclink_reg[128]_net_1 , \mdiclink_reg[127]_net_1 , 
        \mdiclink_reg[126]_net_1 , \mdiclink_reg[125]_net_1 , 
        \mdiclink_reg[124]_net_1 , \mdiclink_reg[123]_net_1 , 
        \mdiclink_reg[122]_net_1 , \mdiclink_reg[121]_net_1 , 
        \mdiclink_reg[120]_net_1 , \mdiclink_reg[119]_net_1 , 
        \mdiclink_reg[118]_net_1 , \mdiclink_reg[117]_net_1 , 
        \mdiclink_reg[116]_net_1 , \mdiclink_reg[115]_net_1 , 
        \mdiclink_reg[114]_net_1 , \mdiclink_reg[113]_net_1 , 
        \mdiclink_reg[112]_net_1 , \mdiclink_reg[111]_net_1 , 
        \mdiclink_reg[110]_net_1 , \mdiclink_reg[109]_net_1 , 
        \mdiclink_reg[108]_net_1 , \mdiclink_reg[107]_net_1 , 
        \mdiclink_reg[106]_net_1 , \mdiclink_reg[105]_net_1 , 
        \mdiclink_reg[104]_net_1 , \mdiclink_reg[103]_net_1 , 
        \mdiclink_reg[102]_net_1 , \mdiclink_reg[101]_net_1 , 
        \mdiclink_reg[100]_net_1 , \mdiclink_reg[99]_net_1 , 
        \mdiclink_reg[98]_net_1 , \mdiclink_reg[97]_net_1 , 
        \mdiclink_reg[96]_net_1 , \mdiclink_reg[95]_net_1 , 
        \mdiclink_reg[94]_net_1 , \mdiclink_reg[93]_net_1 , 
        \mdiclink_reg[92]_net_1 , \mdiclink_reg[91]_net_1 , 
        \mdiclink_reg[90]_net_1 , \mdiclink_reg[89]_net_1 , 
        \mdiclink_reg[88]_net_1 , \mdiclink_reg[87]_net_1 , 
        \mdiclink_reg[86]_net_1 , \mdiclink_reg[85]_net_1 , 
        \mdiclink_reg[84]_net_1 , \mdiclink_reg[83]_net_1 , 
        \mdiclink_reg[82]_net_1 , \mdiclink_reg[81]_net_1 , 
        \mdiclink_reg[80]_net_1 , \mdiclink_reg[79]_net_1 , 
        \mdiclink_reg[78]_net_1 , \mdiclink_reg[77]_net_1 , 
        \mdiclink_reg[76]_net_1 , \mdiclink_reg[75]_net_1 , 
        \mdiclink_reg[74]_net_1 , \mdiclink_reg[73]_net_1 , 
        \mdiclink_reg[72]_net_1 , \mdiclink_reg[71]_net_1 , 
        \mdiclink_reg[70]_net_1 , \mdiclink_reg[69]_net_1 , 
        \mdiclink_reg[68]_net_1 , \mdiclink_reg[67]_net_1 , 
        \mdiclink_reg[66]_net_1 , \mdiclink_reg[65]_net_1 , 
        \mdiclink_reg[64]_net_1 , \mdiclink_reg[63]_net_1 , 
        \mdiclink_reg[62]_net_1 , \mdiclink_reg[61]_net_1 , 
        \mdiclink_reg[60]_net_1 , \mdiclink_reg[59]_net_1 , 
        \mdiclink_reg[58]_net_1 , \mdiclink_reg[57]_net_1 , 
        \mdiclink_reg[56]_net_1 , \mdiclink_reg[55]_net_1 , 
        \mdiclink_reg[54]_net_1 , \mdiclink_reg[53]_net_1 , 
        \mdiclink_reg[52]_net_1 , \mdiclink_reg[51]_net_1 , 
        \mdiclink_reg[50]_net_1 , \mdiclink_reg[49]_net_1 , 
        \mdiclink_reg[48]_net_1 , \mdiclink_reg[47]_net_1 , 
        \mdiclink_reg[46]_net_1 , \mdiclink_reg[45]_net_1 , 
        \mdiclink_reg[44]_net_1 , \mdiclink_reg[43]_net_1 , 
        \mdiclink_reg[42]_net_1 , \mdiclink_reg[41]_net_1 , 
        \mdiclink_reg[40]_net_1 , \mdiclink_reg[39]_net_1 , 
        \mdiclink_reg[38]_net_1 , \mdiclink_reg[37]_net_1 , 
        \mdiclink_reg[36]_net_1 , \mdiclink_reg[35]_net_1 , 
        \mdiclink_reg[34]_net_1 , \mdiclink_reg[33]_net_1 , 
        \mdiclink_reg[32]_net_1 , \mdiclink_reg[31]_net_1 , 
        \mdiclink_reg[30]_net_1 , \mdiclink_reg[29]_net_1 , 
        \mdiclink_reg[28]_net_1 , \mdiclink_reg[27]_net_1 , 
        \mdiclink_reg[26]_net_1 , \mdiclink_reg[25]_net_1 , 
        \mdiclink_reg[24]_net_1 , \mdiclink_reg[23]_net_1 , 
        \mdiclink_reg[22]_net_1 , \mdiclink_reg[21]_net_1 , 
        \mdiclink_reg[20]_net_1 , \mdiclink_reg[19]_net_1 , 
        \mdiclink_reg[18]_net_1 , \mdiclink_reg[17]_net_1 , 
        \mdiclink_reg[16]_net_1 , \mdiclink_reg[15]_net_1 , 
        \mdiclink_reg[14]_net_1 , \mdiclink_reg[13]_net_1 , 
        \mdiclink_reg[12]_net_1 , \mdiclink_reg[11]_net_1 , 
        \mdiclink_reg[10]_net_1 , \mdiclink_reg[9]_net_1 , 
        \mdiclink_reg[8]_net_1 , \mdiclink_reg[7]_net_1 , 
        \mdiclink_reg[6]_net_1 , \mdiclink_reg[5]_net_1 , 
        \mdiclink_reg[4]_net_1 , \mdiclink_reg[3]_net_1 , 
        \mdiclink_reg[2]_net_1 , \mdiclink_reg[1]_net_1 , 
        \mdiclink_reg[0]_net_1 }), .b6_Ocm0rW_0_0_o2({
        \b6_Ocm0rW_0_0_o2[2] }), .b13_nAzGfFM_sLsv3({
        \b13_nAzGfFM_sLsv3[1] }), .IICE_comm2iice_11(
        IICE_comm2iice[11]), .IICE_comm2iice_10(IICE_comm2iice[10]), 
        .IICE_comm2iice_5(IICE_comm2iice[5]), .IICE_comm2iice_0(
        IICE_comm2iice[0]), .IICE_comm2iice_4(IICE_comm2iice[4]), 
        .IICE_comm2iice_9(IICE_comm2iice[9]), .IICE_comm2iice_1(
        IICE_comm2iice[1]), .IICE_comm2iice_3(IICE_comm2iice[3]), 
        .IICE_comm2iice_2(IICE_comm2iice[2]), .IICE_comm2iice_6(
        IICE_comm2iice[6]), .BW_clk_c(BW_clk_c), .b11_PSyil9s_FMZ(
        b11_PSyil9s_FMZ), .b8_SoWGfWYY_i(b8_SoWGfWYY_i), .b8_SoWGfWYY(
        b8_SoWGfWYY), .b10_OFWNT9khFt(b10_OFWNT9khFt), .b7_yYh03wy(
        b7_yYh03wy), .b9_OFWNT9Mxf(b9_OFWNT9Mxf));
    SLE \mdiclink_reg[91]  (.D(\data_from_adc[5] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[91]_net_1 ));
    SLE \mdiclink_reg[352]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[352]_net_1 ));
    SLE \mdiclink_reg[111]  (.D(\data_from_adc[3] [10]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[111]_net_1 ));
    SLE \mdiclink_reg[147]  (.D(\data_from_adc[0] [10]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[147]_net_1 ));
    SLE \mdiclink_reg[34]  (.D(dac1_db_c[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[34]_net_1 ));
    SLE \mdiclink_reg[252]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[252]_net_1 ));
    SLE \mdiclink_reg[198]  (.D(fpga_shift_2[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[198]_net_1 ));
    SLE \mdiclink_reg[146]  (.D(\data_from_adc[0] [11]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[146]_net_1 ));
    SLE \mdiclink_reg[140]  (.D(\data_from_adc[1] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[140]_net_1 ));
    b3_uKr_x b8_uKr_IFLY (.b13_nvmFL_fx2rbuQ({IICE_comm2iice[0], 
        IICE_comm2iice[1], IICE_comm2iice[2], IICE_comm2iice[3], 
        IICE_comm2iice[4], IICE_comm2iice[5]}), .b11_uRrc_9urXBb(
        IICE_comm2iice[6]), .b3_PLy(IICE_comm2iice[7]), .b3_PLF(
        IICE_iice2comm), .b7_PLy_PlM(b4_PLyF), .b12_PSyiBgfDb_bd(
        b8_PSyiBgYG), .b12_PSyi2XfYF_bd(b8_PSyi2XYG), 
        .b14_OFWNT9khWqH_3i(b10_OFWNT9khFt), .b13_PSyiBgfDb_Z4D(
        b7_PSyi3wy), .b13_PSyi2XfYF_Z4D(GND_net_1), 
        .b15_OFWNT9khWqH_R9k(b9_OFWNT9Mxf), .b7_yYh03wy(b7_yYh03wy), 
        .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), .b11_uRrc2XfY_XH(
        b11_uRrc2XfY_XH), .b13_nUTQBgfDb_Z4D(b13_nUTQBgfDb_Z4D), 
        .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), 
        .b16_nYhI39swMeEd_A78(b16_nYhI39swMeEd_A78), .b11_vABZ3qsY_XH(
        b11_vABZ3qsY_XH), .b12_vABZ3qsY_Lyh(b12_vABZ3qsY_Lyh), 
        .b12_ibScJX_E2_bd(b12_ibScJX_E2_bd), .b13_ibScJX_E2_Z4D(
        GND_net_1), .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh));
    SLE \mdiclink_reg[318]  (.D(temp_count[19]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[318]_net_1 ));
    SLE \mdiclink_reg[298]  (.D(temp3[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[298]_net_1 ));
    SLE \mdiclink_reg[294]  (.D(temp3[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[294]_net_1 ));
    SLE \mdiclink_reg[167]  (.D(dds_sin[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[167]_net_1 ));
    SLE \mdiclink_reg[349]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[349]_net_1 ));
    SLE \mdiclink_reg[257]  (.D(temp1[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[257]_net_1 ));
    SLE \mdiclink_reg[166]  (.D(dds_sin[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[166]_net_1 ));
    SLE \mdiclink_reg[1]  (.D(BW_c[13]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[1]_net_1 ));
    SLE \mdiclink_reg[160]  (.D(dds_cos[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[160]_net_1 ));
    SLE \mdiclink_reg[246]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[246]_net_1 ));
    SLE \mdiclink_reg[93]  (.D(\data_from_adc[5] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[93]_net_1 ));
    SLE \mdiclink_reg[69]  (.D(\data_from_adc[7] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[69]_net_1 ));
    SLE \mdiclink_reg[104]  (.D(\data_from_adc[4] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[104]_net_1 ));
    SLE \mdiclink_reg[293]  (.D(temp3[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[293]_net_1 ));
    SLE \mdiclink_reg[112]  (.D(\data_from_adc[3] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[112]_net_1 ));
    SLE \mdiclink_reg[369]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[369]_net_1 ));
    SLE \mdiclink_reg[305]  (.D(temp3_csn_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[305]_net_1 ));
    SLE \mdiclink_reg[179]  (.D(fpga_count[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[179]_net_1 ));
    SLE \mdiclink_reg[340]  (.D(temp_count_data[2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[340]_net_1 ));
    SLE \mdiclink_reg[266]  (.D(temp1[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[266]_net_1 ));
    SLE \mdiclink_reg[229]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[229]_net_1 ));
    SLE \mdiclink_reg[22]  (.D(BW_out_c[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[22]_net_1 ));
    SLE \mdiclink_reg[98]  (.D(\data_from_adc[4] [11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[98]_net_1 ));
    SLE \mdiclink_reg[316]  (.D(temp_count[21]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[316]_net_1 ));
    SLE \mdiclink_reg[201]  (.D(fpga_shift_2[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[201]_net_1 ));
    SLE \mdiclink_reg[188]  (.D(fpga_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[188]_net_1 ));
    SLE \mdiclink_reg[360]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[360]_net_1 ));
    SLE \mdiclink_reg[81]  (.D(\data_from_adc[6] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[81]_net_1 ));
    SLE \mdiclink_reg[288]  (.D(temp2_csn_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[288]_net_1 ));
    SLE \mdiclink_reg[284]  (.D(temp2[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[284]_net_1 ));
    SLE \mdiclink_reg[121]  (.D(\data_from_adc[3] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[121]_net_1 ));
    SLE \mdiclink_reg[96]  (.D(\data_from_adc[5] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[96]_net_1 ));
    SLE \mdiclink_reg[301]  (.D(temp3[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[301]_net_1 ));
    SLE \mdiclink_reg[177]  (.D(fpga_count[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[177]_net_1 ));
    SLE \mdiclink_reg[138]  (.D(\data_from_adc[1] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[138]_net_1 ));
    SLE \mdiclink_reg[210]  (.D(fr_adc_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[210]_net_1 ));
    SLE \mdiclink_reg[176]  (.D(fpga_count[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[176]_net_1 ));
    SLE \mdiclink_reg[283]  (.D(temp2[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[283]_net_1 ));
    SLE \mdiclink_reg[238]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[238]_net_1 ));
    SLE \mdiclink_reg[170]  (.D(dds_sin[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[170]_net_1 ));
    SLE \mdiclink_reg[234]  (.D(freq_11), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[234]_net_1 ));
    SLE \mdiclink_reg[65]  (.D(\data_from_adc[7] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[65]_net_1 ));
    SLE \mdiclink_reg[328]  (.D(temp_count[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[328]_net_1 ));
    SLE \mdiclink_reg[24]  (.D(BW_out_c[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[24]_net_1 ));
    SLE \mdiclink_reg[193]  (.D(fpga_shift_2[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[193]_net_1 ));
    SLE \mdiclink_reg[276]  (.D(temp2[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[276]_net_1 ));
    SLE \mdiclink_reg[39]  (.D(dac1_db_c[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[39]_net_1 ));
    SLE \mdiclink_reg[343]  (.D(temp_sck_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[343]_net_1 ));
    SLE \mdiclink_reg[233]  (.D(VCC_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[233]_net_1 ));
    SLE \mdiclink_reg[83]  (.D(\data_from_adc[6] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[83]_net_1 ));
    SLE \mdiclink_reg[259]  (.D(temp1[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[259]_net_1 ));
    SLE \mdiclink_reg[12]  (.D(BW_c[2]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[12]_net_1 ));
    SLE \mdiclink_reg[122]  (.D(\data_from_adc[2] [11]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[122]_net_1 ));
    SLE \mdiclink_reg[370]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[370]_net_1 ));
    SLE \mdiclink_reg[363]  (.D(freq_6), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[363]_net_1 ));
    SLE \mdiclink_reg[302]  (.D(temp3[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[302]_net_1 ));
    SLE \mdiclink_reg[60]  (.D(\data_from_adc[8] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[60]_net_1 ));
    SLE \mdiclink_reg[334]  (.D(temp_count[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[334]_net_1 ));
    SLE \mdiclink_reg[41]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[41]_net_1 ));
    SLE \mdiclink_reg[215]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[215]_net_1 ));
    SLE \mdiclink_reg[151]  (.D(\data_from_adc[0] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[151]_net_1 ));
    SLE \mdiclink_reg[326]  (.D(temp_count[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[326]_net_1 ));
    SLE \mdiclink_reg[67]  (.D(\data_from_adc[7] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[67]_net_1 ));
    SLE \mdiclink_reg[88]  (.D(\data_from_adc[5] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[88]_net_1 ));
    SLE \mdiclink_reg[202]  (.D(fpga_shift_2[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[202]_net_1 ));
    SLE \mdiclink_reg[195]  (.D(fpga_shift_2[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[195]_net_1 ));
    SLE \mdiclink_reg[4]  (.D(BW_c[10]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[4]_net_1 ));
    SLE \mdiclink_reg[183]  (.D(fpga_count[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[183]_net_1 ));
    SLE \mdiclink_reg[72]  (.D(\data_from_adc[7] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[72]_net_1 ));
    SLE \mdiclink_reg[86]  (.D(\data_from_adc[5] [11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[86]_net_1 ));
    SLE \mdiclink_reg[358]  (.D(freq_11), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[358]_net_1 ));
    SLE \mdiclink_reg[14]  (.D(BW_c[0]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[14]_net_1 ));
    SLE \mdiclink_reg[220]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[220]_net_1 ));
    SLE \mdiclink_reg[207]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[207]_net_1 ));
    SLE \mdiclink_reg[35]  (.D(dac1_db_c[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[35]_net_1 ));
    SLE \mdiclink_reg[133]  (.D(\data_from_adc[2] [0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[133]_net_1 ));
    SLE \mdiclink_reg[43]  (.D(dac_count[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[43]_net_1 ));
    SLE \mdiclink_reg[152]  (.D(\data_from_adc[0] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[152]_net_1 ));
    SLE \mdiclink_reg[144]  (.D(\data_from_adc[1] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[144]_net_1 ));
    SLE \mdiclink_reg[373]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[373]_net_1 ));
    SLE \mdiclink_reg[345]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[345]_net_1 ));
    SLE \mdiclink_reg[74]  (.D(\data_from_adc[6] [11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[74]_net_1 ));
    SLE \mdiclink_reg[164]  (.D(dds_cos[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[164]_net_1 ));
    SLE \mdiclink_reg[356]  (.D(freq_13), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[356]_net_1 ));
    SLE \mdiclink_reg[185]  (.D(fpga_count[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[185]_net_1 ));
    SLE \mdiclink_reg[29]  (.D(BW_out_c[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[29]_net_1 ));
    SLE \mdiclink_reg[365]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[365]_net_1 ));
    SLE \mdiclink_reg[30]  (.D(dac1_clk_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[30]_net_1 ));
    SLE \mdiclink_reg[48]  (.D(dac_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[48]_net_1 ));
    SLE \mdiclink_reg[241]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[241]_net_1 ));
    SLE \mdiclink_reg[225]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[225]_net_1 ));
    SLE \mdiclink_reg[37]  (.D(dac1_db_c[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[37]_net_1 ));
    SLE \mdiclink_reg[46]  (.D(dac_count[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[46]_net_1 ));
    SLE \mdiclink_reg[135]  (.D(\data_from_adc[1] [10]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[135]_net_1 ));
    SLE \mdiclink_reg[261]  (.D(temp1[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[261]_net_1 ));
    SLE \mdiclink_reg[199]  (.D(fpga_shift_2[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[199]_net_1 ));
    SLE \mdiclink_reg[250]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[250]_net_1 ));
    SLE \mdiclink_reg[341]  (.D(temp_count_data[1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[341]_net_1 ));
    SLE \mdiclink_reg[118]  (.D(\data_from_adc[3] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[118]_net_1 ));
    SLE \mdiclink_reg[5]  (.D(BW_c[9]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[5]_net_1 ));
    SLE \mdiclink_reg[218]  (.D(fr_adc_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[218]_net_1 ));
    SLE \mdiclink_reg[214]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[214]_net_1 ));
    SLE \mdiclink_reg[361]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[361]_net_1 ));
    SLE \mdiclink_reg[209]  (.D(fr_adc_count[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[209]_net_1 ));
    SLE \mdiclink_reg[19]  (.D(BW_out_c[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[19]_net_1 ));
    SLE \mdiclink_reg[174]  (.D(temp_sck_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[174]_net_1 ));
    SLE \mdiclink_reg[92]  (.D(\data_from_adc[5] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[92]_net_1 ));
    SLE \mdiclink_reg[25]  (.D(BW_out_c[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[25]_net_1 ));
    SLE \mdiclink_reg[213]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[213]_net_1 ));
    SLE \mdiclink_reg[197]  (.D(fpga_shift_2[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[197]_net_1 ));
    SLE \mdiclink_reg[375]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[375]_net_1 ));
    SLE \mdiclink_reg[3]  (.D(BW_c[11]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[3]_net_1 ));
    SLE \mdiclink_reg[196]  (.D(fpga_shift_2[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[196]_net_1 ));
    SLE \mdiclink_reg[190]  (.D(fpga_shift_2[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[190]_net_1 ));
    SLE \mdiclink_reg[342]  (.D(temp_count_data[0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[342]_net_1 ));
    SLE \mdiclink_reg[255]  (.D(temp1[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[255]_net_1 ));
    SLE \mdiclink_reg[101]  (.D(\data_from_adc[4] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[101]_net_1 ));
    SLE \mdiclink_reg[189]  (.D(fpga_count[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[189]_net_1 ));
    SLE \mdiclink_reg[337]  (.D(temp_count[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[337]_net_1 ));
    SLE \mdiclink_reg[314]  (.D(temp_count[23]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[314]_net_1 ));
    SLE \mdiclink_reg[271]  (.D(temp1_csn_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[271]_net_1 ));
    SLE \mdiclink_reg[362]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[362]_net_1 ));
    SLE \mdiclink_reg[296]  (.D(temp3[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[296]_net_1 ));
    SLE \mdiclink_reg[242]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[242]_net_1 ));
    SLE \mdiclink_reg[308]  (.D(temp_count[29]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[308]_net_1 ));
    SLE \mdiclink_reg[139]  (.D(\data_from_adc[1] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[139]_net_1 ));
    SLE \mdiclink_reg[79]  (.D(\data_from_adc[6] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[79]_net_1 ));
    SLE \mdiclink_reg[20]  (.D(BW_out_c[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[20]_net_1 ));
    SLE \mdiclink_reg[94]  (.D(\data_from_adc[5] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[94]_net_1 ));
    SLE \mdiclink_reg[371]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[371]_net_1 ));
    SLE \mdiclink_reg[27]  (.D(BW_out_c[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[27]_net_1 ));
    SLE \mdiclink_reg[262]  (.D(temp1[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[262]_net_1 ));
    SLE \mdiclink_reg[247]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[247]_net_1 ));
    SLE \mdiclink_reg[128]  (.D(\data_from_adc[2] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[128]_net_1 ));
    SLE \mdiclink_reg[51]  (.D(\data_from_adc[8] [10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[51]_net_1 ));
    SLE \mdiclink_reg[187]  (.D(fpga_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[187]_net_1 ));
    SLE \mdiclink_reg[228]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[228]_net_1 ));
    SLE \mdiclink_reg[15]  (.D(BW_out_c[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[15]_net_1 ));
    SLE \mdiclink_reg[102]  (.D(\data_from_adc[4] [7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[102]_net_1 ));
    SLE \mdiclink_reg[224]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[224]_net_1 ));
    SLE \mdiclink_reg[186]  (.D(fpga_count[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[186]_net_1 ));
    SLE \mdiclink_reg[180]  (.D(fpga_count[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[180]_net_1 ));
    SLE \mdiclink_reg[113]  (.D(\data_from_adc[3] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[113]_net_1 ));
    SLE \mdiclink_reg[267]  (.D(temp1[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[267]_net_1 ));
    SLE \mdiclink_reg[137]  (.D(\data_from_adc[1] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[137]_net_1 ));
    SLE \mdiclink_reg[306]  (.D(temp_count[31]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[306]_net_1 ));
    SLE \mdiclink_reg[223]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[223]_net_1 ));
    SLE \mdiclink_reg[286]  (.D(temp2[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[286]_net_1 ));
    SLE \mdiclink_reg[136]  (.D(\data_from_adc[1] [9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[136]_net_1 ));
    SLE \mdiclink_reg[82]  (.D(\data_from_adc[6] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[82]_net_1 ));
    SLE \mdiclink_reg[130]  (.D(\data_from_adc[2] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[130]_net_1 ));
    SLE \mdiclink_reg[372]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[372]_net_1 ));
    SLE \mdiclink_reg[10]  (.D(BW_c[4]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[10]_net_1 ));
    SLE \mdiclink_reg[75]  (.D(\data_from_adc[6] [10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[75]_net_1 ));
    SLE \mdiclink_reg[339]  (.D(temp_count_data[3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[339]_net_1 ));
    SLE \mdiclink_reg[0]  (.D(BW_c[14]), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[0]_net_1 ));
    SLE \mdiclink_reg[324]  (.D(temp_count[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[324]_net_1 ));
    SLE \mdiclink_reg[53]  (.D(\data_from_adc[8] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[53]_net_1 ));
    SLE \mdiclink_reg[236]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[236]_net_1 ));
    SLE \mdiclink_reg[200]  (.D(fpga_shift_2[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[200]_net_1 ));
    SLE \mdiclink_reg[17]  (.D(BW_out_c[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[17]_net_1 ));
    SLE \mdiclink_reg[272]  (.D(temp2[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[272]_net_1 ));
    SLE \mdiclink_reg[158]  (.D(dds_cos[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[158]_net_1 ));
    SLE \mdiclink_reg[115]  (.D(\data_from_adc[3] [6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[115]_net_1 ));
    SLE \mdiclink_reg[330]  (.D(temp_count[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[330]_net_1 ));
    SLE \mdiclink_reg[258]  (.D(temp1[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[258]_net_1 ));
    SLE \mdiclink_reg[254]  (.D(sdv_count[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[254]_net_1 ));
    SLE \mdiclink_reg[84]  (.D(\data_from_adc[6] [1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[84]_net_1 ));
    SLE \mdiclink_reg[277]  (.D(temp2[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[277]_net_1 ));
    SLE \mdiclink_reg[58]  (.D(\data_from_adc[8] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[58]_net_1 ));
    SLE \mdiclink_reg[70]  (.D(\data_from_adc[7] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[70]_net_1 ));
    SLE \mdiclink_reg[249]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[249]_net_1 ));
    SLE \mdiclink_reg[253]  (.D(sdv_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[253]_net_1 ));
    SLE \mdiclink_reg[123]  (.D(\data_from_adc[2] [10]), .CLK(BW_clk_c)
        , .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[123]_net_1 ));
    SLE \mdiclink_reg[77]  (.D(\data_from_adc[6] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[77]_net_1 ));
    SLE \mdiclink_reg[56]  (.D(\data_from_adc[8] [5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[56]_net_1 ));
    SLE \mdiclink_reg[99]  (.D(\data_from_adc[4] [10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[99]_net_1 ));
    SLE \mdiclink_reg[42]  (.D(dac_count[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[42]_net_1 ));
    SLE \mdiclink_reg[205]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[205]_net_1 ));
    SLE \mdiclink_reg[269]  (.D(temp1[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[269]_net_1 ));
    SLE \mdiclink_reg[141]  (.D(\data_from_adc[1] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[141]_net_1 ));
    SLE \mdiclink_reg[354]  (.D(freq_15), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[354]_net_1 ));
    SLE \mdiclink_reg[7]  (.D(BW_c[7]), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[7]_net_1 ));
    SLE \mdiclink_reg[317]  (.D(temp_count[20]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[317]_net_1 ));
    SLE \mdiclink_reg[161]  (.D(dds_cos[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[161]_net_1 ));
    SLE \mdiclink_reg[348]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[348]_net_1 ));
    SLE \mdiclink_reg[333]  (.D(temp_count[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[333]_net_1 ));
    SLE \mdiclink_reg[194]  (.D(fpga_shift_2[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[194]_net_1 ));
    SLE \mdiclink_reg[119]  (.D(\data_from_adc[3] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[119]_net_1 ));
    SLE \mdiclink_reg[44]  (.D(dac_count[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[44]_net_1 ));
    SLE \mdiclink_reg[125]  (.D(\data_from_adc[2] [8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[125]_net_1 ));
    SLE \mdiclink_reg[368]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[368]_net_1 ));
    SLE \mdiclink_reg[95]  (.D(\data_from_adc[5] [2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[95]_net_1 ));
    SLE \mdiclink_reg[153]  (.D(\data_from_adc[0] [4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[153]_net_1 ));
    SLE \mdiclink_reg[142]  (.D(\data_from_adc[1] [3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[142]_net_1 ));
    
endmodule


module b9_ORbIwXaEF_32s_2494704002_0s_x_0(
       b3_ORb_0,
       tck,
       b6_nv_0CC,
       b10_nv_ywKMm9X,
       b12_ORbIwXaEF_bd,
       b8_nv_ZmCtY
    );
output b3_ORb_0;
input  tck;
input  b6_nv_0CC;
input  b10_nv_ywKMm9X;
input  b12_ORbIwXaEF_bd;
input  b8_nv_ZmCtY;

    wire b3_ORb_7_net_1, N_458_i, \b3_ORb[23]_net_1 , VCC_net_1, 
        \b3_ORb[24]_net_1 , \b3_ORb_or[7]_net_1 , GND_net_1, 
        \b3_ORb[25]_net_1 , \b3_ORb[26]_net_1 , \b3_ORb[27]_net_1 , 
        \b3_ORb[28]_net_1 , \b3_ORb[29]_net_1 , \b3_ORb[30]_net_1 , 
        \b3_ORb[31]_net_1 , \b3_ORb[32]_net_1 , \b3_ORb[8]_net_1 , 
        \b3_ORb[9]_net_1 , \b3_ORb[10]_net_1 , \b3_ORb[11]_net_1 , 
        \b3_ORb[12]_net_1 , \b3_ORb[13]_net_1 , \b3_ORb[14]_net_1 , 
        \b3_ORb[15]_net_1 , \b3_ORb[16]_net_1 , \b3_ORb[17]_net_1 , 
        \b3_ORb[18]_net_1 , \b3_ORb[19]_net_1 , \b3_ORb[20]_net_1 , 
        \b3_ORb[21]_net_1 , \b3_ORb[22]_net_1 , \b3_ORb[2]_net_1 , 
        \b3_ORb[3]_net_1 , \b3_ORb[4]_net_1 , \b3_ORb[5]_net_1 , 
        \b3_ORb[6]_net_1 , \b3_ORb[7]_net_1 , un1_b3_ORb9_i_0;
    
    SLE \b3_ORb[7]  (.D(\b3_ORb[8]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[7]_net_1 ));
    SLE \b3_ORb[9]  (.D(\b3_ORb[10]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[9]_net_1 ));
    SLE \b3_ORb[3]  (.D(\b3_ORb[4]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[3]_net_1 ));
    SLE \b3_ORb[23]  (.D(\b3_ORb[24]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[23]_net_1 ));
    SLE \b3_ORb[22]  (.D(\b3_ORb[23]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[22]_net_1 ));
    SLE \b3_ORb[1]  (.D(\b3_ORb[2]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(b3_ORb_0));
    SLE \b3_ORb[10]  (.D(\b3_ORb[11]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[10]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_458_i_0 (.A(b3_ORb_7_net_1), .Y(N_458_i));
    CFG2 #( .INIT(4'hE) )  \b3_ORb_or[7]  (.A(b3_ORb_7_net_1), .B(
        un1_b3_ORb9_i_0), .Y(\b3_ORb_or[7]_net_1 ));
    SLE \b3_ORb[16]  (.D(\b3_ORb[17]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[16]_net_1 ));
    SLE \b3_ORb[11]  (.D(\b3_ORb[12]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[11]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  b3_ORb_7 (.A(b10_nv_ywKMm9X), .B(
        b12_ORbIwXaEF_bd), .Y(b3_ORb_7_net_1));
    SLE \b3_ORb[17]  (.D(\b3_ORb[18]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[17]_net_1 ));
    SLE \b3_ORb[5]  (.D(\b3_ORb[6]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[5]_net_1 ));
    SLE \b3_ORb[28]  (.D(\b3_ORb[29]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[28]_net_1 ));
    SLE \b3_ORb[6]  (.D(\b3_ORb[7]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[6]_net_1 ));
    SLE \b3_ORb[29]  (.D(\b3_ORb[30]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[29]_net_1 ));
    SLE \b3_ORb[13]  (.D(\b3_ORb[14]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[13]_net_1 ));
    SLE \b3_ORb[12]  (.D(\b3_ORb[13]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[12]_net_1 ));
    SLE \b3_ORb[24]  (.D(\b3_ORb[25]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[24]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hC8) )  un1_b3_ORb9_i (.A(b10_nv_ywKMm9X), .B(
        b12_ORbIwXaEF_bd), .C(b8_nv_ZmCtY), .Y(un1_b3_ORb9_i_0));
    SLE \b3_ORb[2]  (.D(\b3_ORb[3]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[2]_net_1 ));
    SLE \b3_ORb[25]  (.D(\b3_ORb[26]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[25]_net_1 ));
    SLE \b3_ORb[30]  (.D(\b3_ORb[31]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[30]_net_1 ));
    SLE \b3_ORb[18]  (.D(\b3_ORb[19]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[18]_net_1 ));
    SLE \b3_ORb[20]  (.D(\b3_ORb[21]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[20]_net_1 ));
    SLE \b3_ORb[19]  (.D(\b3_ORb[20]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[19]_net_1 ));
    SLE \b3_ORb[31]  (.D(\b3_ORb[32]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[31]_net_1 ));
    SLE \b3_ORb[14]  (.D(\b3_ORb[15]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[14]_net_1 ));
    SLE \b3_ORb[26]  (.D(\b3_ORb[27]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[26]_net_1 ));
    SLE \b3_ORb[4]  (.D(\b3_ORb[5]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[4]_net_1 ));
    SLE \b3_ORb[21]  (.D(\b3_ORb[22]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[21]_net_1 ));
    SLE \b3_ORb[8]  (.D(\b3_ORb[9]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[8]_net_1 ));
    SLE \b3_ORb[15]  (.D(\b3_ORb[16]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[15]_net_1 ));
    SLE \b3_ORb[27]  (.D(\b3_ORb[28]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[27]_net_1 ));
    SLE \b3_ORb[32]  (.D(b6_nv_0CC), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[32]_net_1 ));
    
endmodule


module jtag_interface_x_0(
       b9_OvyH3_saL,
       b11_uRrc_WYOFjZ,
       b11_uRrc_9urXBb,
       dr2_tck_i,
       tdo_sig,
       b12_ORbIwXaEF_bd,
       IICE_iice2comm,
       b10_8Kz_fFfsjX,
       b5_OvyH3,
       b8_nv_ZmCtY,
       b7_nFG0rDY,
       b10_nv_ywKMm9X,
       hcr_update,
       ch_update,
       b6_nv_0CC,
       atrstb,
       atdo,
       atdi,
       atms,
       atck
    );
input  [0:0] b9_OvyH3_saL;
input  [0:0] b11_uRrc_WYOFjZ;
output [0:0] b11_uRrc_9urXBb;
output dr2_tck_i;
input  tdo_sig;
input  b12_ORbIwXaEF_bd;
input  IICE_iice2comm;
output b10_8Kz_fFfsjX;
output b5_OvyH3;
output b8_nv_ZmCtY;
output b7_nFG0rDY;
output b10_nv_ywKMm9X;
output hcr_update;
output ch_update;
output b6_nv_0CC;
input  atrstb;
output atdo;
input  atdi;
input  atms;
input  atck;

    wire identify_clk_int, b3_1Um, b9_96_cLqgOF4_net_1, 
        b9_PLF_6lNa2_1_net_1, b9_PLF_6lNa2_net_1, b9_96_cLqgOF3_net_1, 
        \b6_uS_MrX[2] , \b6_uS_MrX[3] , b9_96_cLqgOF4_2, 
        \b6_uS_MrX[0] , \b6_uS_MrX[4] , \b6_uS_MrX[1] , 
        identify_clk2_no_clk_buffer_needed, \UIREGdummy[0] , 
        \UIREGdummy[7] , URSTBdummy, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h0008) )  b9_96_cLqgOF3 (.A(\b6_uS_MrX[0] ), .B(
        b9_96_cLqgOF4_2), .C(\b6_uS_MrX[4] ), .D(\b6_uS_MrX[1] ), .Y(
        b9_96_cLqgOF3_net_1));
    CFG2 #( .INIT(4'h8) )  b10_8Kz_fFfsjX_inst_1 (.A(
        b9_96_cLqgOF4_net_1), .B(b3_1Um), .Y(b10_8Kz_fFfsjX));
    CFG3 #( .INIT(8'h80) )  b10_nv_ywKMm9X_inst_1 (.A(b3_1Um), .B(
        b9_96_cLqgOF3_net_1), .C(b7_nFG0rDY), .Y(b10_nv_ywKMm9X));
    GND GND (.Y(GND_net_1));
    UJTAG b9_Rcmi_KsDw (.UDRCAP(b7_nFG0rDY), .UDRSH(b5_OvyH3), .UDRUPD(
        identify_clk2_no_clk_buffer_needed), .UIREG({\UIREGdummy[7] , 
        b3_1Um, \b6_uS_MrX[4] , \b6_uS_MrX[3] , \b6_uS_MrX[2] , 
        \b6_uS_MrX[1] , \b6_uS_MrX[0] , \UIREGdummy[0] }), .URSTB(
        URSTBdummy), .UDRCK(identify_clk_int), .UTDI(b6_nv_0CC), .UTDO(
        b9_PLF_6lNa2_net_1), .TDI(atdi), .TMS(atms), .TCK(atck), 
        .TRSTB(atrstb), .TDO(atdo));
    CFG3 #( .INIT(8'h80) )  b8_nv_ZmCtY_inst_1 (.A(b3_1Um), .B(
        b9_96_cLqgOF3_net_1), .C(b5_OvyH3), .Y(b8_nv_ZmCtY));
    CFG3 #( .INIT(8'h80) )  b9_nv_oQwfYF_3 (.A(
        identify_clk2_no_clk_buffer_needed), .B(b9_96_cLqgOF3_net_1), 
        .C(b3_1Um), .Y(ch_update));
    CFG2 #( .INIT(4'h8) )  b10_8Kz_rKlrtX_3 (.A(b10_8Kz_fFfsjX), .B(
        identify_clk2_no_clk_buffer_needed), .Y(hcr_update));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h4F7F) )  b9_PLF_6lNa2_1 (.A(tdo_sig), .B(
        b12_ORbIwXaEF_bd), .C(b9_96_cLqgOF3_net_1), .D(IICE_iice2comm), 
        .Y(b9_PLF_6lNa2_1_net_1));
    CFG2 #( .INIT(4'h1) )  b9_96_cLqgOF3_2 (.A(\b6_uS_MrX[2] ), .B(
        \b6_uS_MrX[3] ), .Y(b9_96_cLqgOF4_2));
    CLKINT jtag_clkint_prim (.A(identify_clk_int), .Y(dr2_tck_i));
    CFG4 #( .INIT(16'h0400) )  b9_96_cLqgOF4 (.A(\b6_uS_MrX[0] ), .B(
        b9_96_cLqgOF4_2), .C(\b6_uS_MrX[4] ), .D(\b6_uS_MrX[1] ), .Y(
        b9_96_cLqgOF4_net_1));
    CFG3 #( .INIT(8'h80) )  \b11_uRrc_9urXBb[0]  (.A(
        b11_uRrc_WYOFjZ[0]), .B(b3_1Um), .C(b9_96_cLqgOF3_net_1), .Y(
        b11_uRrc_9urXBb[0]));
    CFG4 #( .INIT(16'h808C) )  b9_PLF_6lNa2 (.A(b9_OvyH3_saL[0]), .B(
        b3_1Um), .C(b9_96_cLqgOF4_net_1), .D(b9_PLF_6lNa2_1_net_1), .Y(
        b9_PLF_6lNa2_net_1));
    
endmodule


module b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0(
       b11_uRrc_WYOFjZ,
       b13_nvmFL_fx2rbuQ,
       b9_OvyH3_saL_0,
       dr2_tck,
       b6_nv_0CC,
       hcr_update,
       b10_8Kz_fFfsjX,
       b12_ORbIwXaEF_bd,
       b7_nFG0rDY,
       b5_OvyH3
    );
output [0:0] b11_uRrc_WYOFjZ;
output [5:0] b13_nvmFL_fx2rbuQ;
output b9_OvyH3_saL_0;
input  dr2_tck;
input  b6_nv_0CC;
input  hcr_update;
input  b10_8Kz_fFfsjX;
output b12_ORbIwXaEF_bd;
input  b7_nFG0rDY;
input  b5_OvyH3;

    wire \b9_OvyH3_saL[1]_net_1 , VCC_net_1, \b9_OvyH3_saL[2]_net_1 , 
        b9_OvyH3_saL_0_sqmuxa_net_1, GND_net_1, 
        \b9_OvyH3_saL[3]_net_1 , \b9_OvyH3_saL[4]_net_1 , 
        \b9_OvyH3_saL[5]_net_1 , \b9_OvyH3_saL[6]_net_1 , 
        \b9_OvyH3_saL[7]_net_1 ;
    
    SLE \genblk1.b10_dZst39_EF3[5]  (.D(\b9_OvyH3_saL[5]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[4]));
    SLE \genblk1.b10_dZst39_EF3[4]  (.D(\b9_OvyH3_saL[4]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[3]));
    SLE \genblk1.b10_dZst39_EF3[3]  (.D(\b9_OvyH3_saL[3]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[2]));
    SLE \genblk1.b10_dZst39_EF3[1]  (.D(\b9_OvyH3_saL[1]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[0]));
    SLE \b9_OvyH3_saL[6]  (.D(\b9_OvyH3_saL[7]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[6]_net_1 ));
    SLE \b9_OvyH3_saL[3]  (.D(\b9_OvyH3_saL[4]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[3]_net_1 ));
    SLE \genblk1.b10_dZst39_EF3[0]  (.D(b9_OvyH3_saL_0), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b11_uRrc_WYOFjZ[0]));
    GND GND (.Y(GND_net_1));
    SLE \genblk1.b10_dZst39_EF3[7]  (.D(\b9_OvyH3_saL[7]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b12_ORbIwXaEF_bd));
    SLE \b9_OvyH3_saL[5]  (.D(\b9_OvyH3_saL[6]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[5]_net_1 ));
    SLE \genblk1.b10_dZst39_EF3[6]  (.D(\b9_OvyH3_saL[6]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[5]));
    SLE \genblk1.b10_dZst39_EF3[2]  (.D(\b9_OvyH3_saL[2]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[1]));
    SLE \b9_OvyH3_saL[7]  (.D(b6_nv_0CC), .CLK(dr2_tck), .EN(
        b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b9_OvyH3_saL[7]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \b9_OvyH3_saL[1]  (.D(\b9_OvyH3_saL[2]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[1]_net_1 ));
    SLE \b9_OvyH3_saL[0]  (.D(\b9_OvyH3_saL[1]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b9_OvyH3_saL_0));
    SLE \b9_OvyH3_saL[4]  (.D(\b9_OvyH3_saL[5]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[4]_net_1 ));
    SLE \b9_OvyH3_saL[2]  (.D(\b9_OvyH3_saL[3]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[2]_net_1 ));
    CFG3 #( .INIT(8'h40) )  b9_OvyH3_saL_0_sqmuxa (.A(b7_nFG0rDY), .B(
        b5_OvyH3), .C(b10_8Kz_fFfsjX), .Y(b9_OvyH3_saL_0_sqmuxa_net_1));
    
endmodule


module comm_block_x(
       IICE_comm2iice,
       IICE_iice2comm,
       atck,
       atdi,
       atdo,
       atms,
       atrstb
    );
output [0:11] IICE_comm2iice;
input  IICE_iice2comm;
input  atck;
input  atdi;
output atdo;
input  atms;
input  atrstb;

    wire hcr_update, b10_8Kz_fFfsjX, \b11_uRrc_WYOFjZ[0] , 
        b12_ORbIwXaEF_bd, tdo_sig, \jtagi.b7_nFG0rDY , 
        \jtagi.b5_OvyH3 , GND_net_1, VCC_net_1, 
        \b7_Rcmi_ql.b9_OvyH3_saL[0] ;
    
    VCC VCC (.Y(VCC_net_1));
    b9_ORbIwXaEF_32s_2494704002_0s_x_0 b9_ORb_xNywD (.b3_ORb_0(tdo_sig)
        , .tck(IICE_comm2iice[11]), .b6_nv_0CC(IICE_comm2iice[7]), 
        .b10_nv_ywKMm9X(IICE_comm2iice[9]), .b12_ORbIwXaEF_bd(
        b12_ORbIwXaEF_bd), .b8_nv_ZmCtY(IICE_comm2iice[10]));
    jtag_interface_x_0 jtagi (.b9_OvyH3_saL({
        \b7_Rcmi_ql.b9_OvyH3_saL[0] }), .b11_uRrc_WYOFjZ({
        \b11_uRrc_WYOFjZ[0] }), .b11_uRrc_9urXBb({IICE_comm2iice[6]}), 
        .dr2_tck_i(IICE_comm2iice[11]), .tdo_sig(tdo_sig), 
        .b12_ORbIwXaEF_bd(b12_ORbIwXaEF_bd), .IICE_iice2comm(
        IICE_iice2comm), .b10_8Kz_fFfsjX(b10_8Kz_fFfsjX), .b5_OvyH3(
        \jtagi.b5_OvyH3 ), .b8_nv_ZmCtY(IICE_comm2iice[10]), 
        .b7_nFG0rDY(\jtagi.b7_nFG0rDY ), .b10_nv_ywKMm9X(
        IICE_comm2iice[9]), .hcr_update(hcr_update), .ch_update(
        IICE_comm2iice[8]), .b6_nv_0CC(IICE_comm2iice[7]), .atrstb(
        atrstb), .atdo(atdo), .atdi(atdi), .atms(atms), .atck(atck));
    GND GND (.Y(GND_net_1));
    b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0 b7_Rcmi_ql 
        (.b11_uRrc_WYOFjZ({\b11_uRrc_WYOFjZ[0] }), .b13_nvmFL_fx2rbuQ({
        IICE_comm2iice[0], IICE_comm2iice[1], IICE_comm2iice[2], 
        IICE_comm2iice[3], IICE_comm2iice[4], IICE_comm2iice[5]}), 
        .b9_OvyH3_saL_0(\b7_Rcmi_ql.b9_OvyH3_saL[0] ), .dr2_tck(
        IICE_comm2iice[11]), .b6_nv_0CC(IICE_comm2iice[7]), 
        .hcr_update(hcr_update), .b10_8Kz_fFfsjX(b10_8Kz_fFfsjX), 
        .b12_ORbIwXaEF_bd(b12_ORbIwXaEF_bd), .b7_nFG0rDY(
        \jtagi.b7_nFG0rDY ), .b5_OvyH3(\jtagi.b5_OvyH3 ));
    
endmodule


module syn_identify_core0_0(
       BW_c,
       BW_out_c,
       dac_count,
       dac1_db_c,
       \data_from_adc[8] ,
       \data_from_adc[7] ,
       \data_from_adc[6] ,
       \data_from_adc[4] ,
       \data_from_adc[5] ,
       \data_from_adc[3] ,
       \data_from_adc[2] ,
       \data_from_adc[1] ,
       \data_from_adc[0] ,
       fpga_count,
       fr_adc_count,
       fpga_shift_2,
       sdv_count,
       temp1,
       temp2,
       temp3,
       temp_count_data,
       temp_count,
       dds_sin,
       dds_cos,
       freq_2,
       freq_14,
       freq_15,
       freq_0,
       freq_1,
       freq_6,
       freq_10,
       freq_11,
       freq_13,
       atck,
       atdi,
       atdo,
       atms,
       atrstb,
       BW_clk_c,
       clk_dac2,
       dac1_clk_c,
       temp_sck_c,
       temp1_csn_c,
       temp2_csn_c,
       temp3_csn_c,
       temp_so_c
    );
input  [14:0] BW_c;
input  [14:0] BW_out_c;
input  [7:1] dac_count;
input  [13:5] dac1_db_c;
input  [11:0] \data_from_adc[8] ;
input  [11:0] \data_from_adc[7] ;
input  [11:0] \data_from_adc[6] ;
input  [11:0] \data_from_adc[4] ;
input  [11:0] \data_from_adc[5] ;
input  [11:0] \data_from_adc[3] ;
input  [11:0] \data_from_adc[2] ;
input  [11:0] \data_from_adc[1] ;
input  [11:0] \data_from_adc[0] ;
input  [14:0] fpga_count;
input  [3:1] fr_adc_count;
input  [14:0] fpga_shift_2;
input  [1:0] sdv_count;
input  [15:0] temp1;
input  [15:0] temp2;
input  [15:0] temp3;
input  [4:0] temp_count_data;
input  [31:0] temp_count;
input  [7:0] dds_sin;
input  [7:0] dds_cos;
input  freq_2;
input  freq_14;
input  freq_15;
input  freq_0;
input  freq_1;
input  freq_6;
input  freq_10;
input  freq_11;
input  freq_13;
input  atck;
input  atdi;
output atdo;
input  atms;
input  atrstb;
input  BW_clk_c;
input  clk_dac2;
input  dac1_clk_c;
input  temp_sck_c;
input  temp1_csn_c;
input  temp2_csn_c;
input  temp3_csn_c;
input  temp_so_c;

    wire \IICE_comm2iice[11] , \IICE_comm2iice[10] , 
        \IICE_comm2iice[9] , \IICE_comm2iice[8] , \IICE_comm2iice[7] , 
        \IICE_comm2iice[6] , \IICE_comm2iice[5] , \IICE_comm2iice[4] , 
        \IICE_comm2iice[3] , \IICE_comm2iice[2] , \IICE_comm2iice[1] , 
        \IICE_comm2iice[0] , IICE_iice2comm, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    IICE_x IICE_INST (.BW_c({BW_c[14], BW_c[13], BW_c[12], BW_c[11], 
        BW_c[10], BW_c[9], BW_c[8], BW_c[7], BW_c[6], BW_c[5], BW_c[4], 
        BW_c[3], BW_c[2], BW_c[1], BW_c[0]}), .BW_out_c({BW_out_c[14], 
        BW_out_c[13], BW_out_c[12], BW_out_c[11], BW_out_c[10], 
        BW_out_c[9], BW_out_c[8], BW_out_c[7], BW_out_c[6], 
        BW_out_c[5], BW_out_c[4], BW_out_c[3], BW_out_c[2], 
        BW_out_c[1], BW_out_c[0]}), .dac_count({dac_count[7], 
        dac_count[6], dac_count[5], dac_count[4], dac_count[3], 
        dac_count[2], dac_count[1]}), .dac1_db_c({dac1_db_c[13], 
        dac1_db_c[12], dac1_db_c[11], dac1_db_c[10], dac1_db_c[9], 
        dac1_db_c[8], dac1_db_c[7], dac1_db_c[6], dac1_db_c[5]}), 
        .\data_from_adc[8] ({\data_from_adc[8] [11], 
        \data_from_adc[8] [10], \data_from_adc[8] [9], 
        \data_from_adc[8] [8], \data_from_adc[8] [7], 
        \data_from_adc[8] [6], \data_from_adc[8] [5], 
        \data_from_adc[8] [4], \data_from_adc[8] [3], 
        \data_from_adc[8] [2], \data_from_adc[8] [1], 
        \data_from_adc[8] [0]}), .\data_from_adc[7] ({
        \data_from_adc[7] [11], \data_from_adc[7] [10], 
        \data_from_adc[7] [9], \data_from_adc[7] [8], 
        \data_from_adc[7] [7], \data_from_adc[7] [6], 
        \data_from_adc[7] [5], \data_from_adc[7] [4], 
        \data_from_adc[7] [3], \data_from_adc[7] [2], 
        \data_from_adc[7] [1], \data_from_adc[7] [0]}), 
        .\data_from_adc[6] ({\data_from_adc[6] [11], 
        \data_from_adc[6] [10], \data_from_adc[6] [9], 
        \data_from_adc[6] [8], \data_from_adc[6] [7], 
        \data_from_adc[6] [6], \data_from_adc[6] [5], 
        \data_from_adc[6] [4], \data_from_adc[6] [3], 
        \data_from_adc[6] [2], \data_from_adc[6] [1], 
        \data_from_adc[6] [0]}), .\data_from_adc[4] ({
        \data_from_adc[4] [11], \data_from_adc[4] [10], 
        \data_from_adc[4] [9], \data_from_adc[4] [8], 
        \data_from_adc[4] [7], \data_from_adc[4] [6], 
        \data_from_adc[4] [5], \data_from_adc[4] [4], 
        \data_from_adc[4] [3], \data_from_adc[4] [2], 
        \data_from_adc[4] [1], \data_from_adc[4] [0]}), 
        .\data_from_adc[5] ({\data_from_adc[5] [11], 
        \data_from_adc[5] [10], \data_from_adc[5] [9], 
        \data_from_adc[5] [8], \data_from_adc[5] [7], 
        \data_from_adc[5] [6], \data_from_adc[5] [5], 
        \data_from_adc[5] [4], \data_from_adc[5] [3], 
        \data_from_adc[5] [2], \data_from_adc[5] [1], 
        \data_from_adc[5] [0]}), .\data_from_adc[3] ({
        \data_from_adc[3] [11], \data_from_adc[3] [10], 
        \data_from_adc[3] [9], \data_from_adc[3] [8], 
        \data_from_adc[3] [7], \data_from_adc[3] [6], 
        \data_from_adc[3] [5], \data_from_adc[3] [4], 
        \data_from_adc[3] [3], \data_from_adc[3] [2], 
        \data_from_adc[3] [1], \data_from_adc[3] [0]}), 
        .\data_from_adc[2] ({\data_from_adc[2] [11], 
        \data_from_adc[2] [10], \data_from_adc[2] [9], 
        \data_from_adc[2] [8], \data_from_adc[2] [7], 
        \data_from_adc[2] [6], \data_from_adc[2] [5], 
        \data_from_adc[2] [4], \data_from_adc[2] [3], 
        \data_from_adc[2] [2], \data_from_adc[2] [1], 
        \data_from_adc[2] [0]}), .\data_from_adc[1] ({
        \data_from_adc[1] [11], \data_from_adc[1] [10], 
        \data_from_adc[1] [9], \data_from_adc[1] [8], 
        \data_from_adc[1] [7], \data_from_adc[1] [6], 
        \data_from_adc[1] [5], \data_from_adc[1] [4], 
        \data_from_adc[1] [3], \data_from_adc[1] [2], 
        \data_from_adc[1] [1], \data_from_adc[1] [0]}), 
        .\data_from_adc[0] ({\data_from_adc[0] [11], 
        \data_from_adc[0] [10], \data_from_adc[0] [9], 
        \data_from_adc[0] [8], \data_from_adc[0] [7], 
        \data_from_adc[0] [6], \data_from_adc[0] [5], 
        \data_from_adc[0] [4], \data_from_adc[0] [3], 
        \data_from_adc[0] [2], \data_from_adc[0] [1], 
        \data_from_adc[0] [0]}), .fpga_count({fpga_count[14], 
        fpga_count[13], fpga_count[12], fpga_count[11], fpga_count[10], 
        fpga_count[9], fpga_count[8], fpga_count[7], fpga_count[6], 
        fpga_count[5], fpga_count[4], fpga_count[3], fpga_count[2], 
        fpga_count[1], fpga_count[0]}), .fr_adc_count({fr_adc_count[3], 
        fr_adc_count[2], fr_adc_count[1]}), .fpga_shift_2({
        fpga_shift_2[14], fpga_shift_2[13], fpga_shift_2[12], 
        fpga_shift_2[11], fpga_shift_2[10], fpga_shift_2[9], 
        fpga_shift_2[8], fpga_shift_2[7], fpga_shift_2[6], 
        fpga_shift_2[5], fpga_shift_2[4], fpga_shift_2[3], 
        fpga_shift_2[2], fpga_shift_2[1], fpga_shift_2[0]}), 
        .sdv_count({sdv_count[1], sdv_count[0]}), .temp1({temp1[15], 
        temp1[14], temp1[13], temp1[12], temp1[11], temp1[10], 
        temp1[9], temp1[8], temp1[7], temp1[6], temp1[5], temp1[4], 
        temp1[3], temp1[2], temp1[1], temp1[0]}), .temp2({temp2[15], 
        temp2[14], temp2[13], temp2[12], temp2[11], temp2[10], 
        temp2[9], temp2[8], temp2[7], temp2[6], temp2[5], temp2[4], 
        temp2[3], temp2[2], temp2[1], temp2[0]}), .temp3({temp3[15], 
        temp3[14], temp3[13], temp3[12], temp3[11], temp3[10], 
        temp3[9], temp3[8], temp3[7], temp3[6], temp3[5], temp3[4], 
        temp3[3], temp3[2], temp3[1], temp3[0]}), .temp_count_data({
        temp_count_data[4], temp_count_data[3], temp_count_data[2], 
        temp_count_data[1], temp_count_data[0]}), .temp_count({
        temp_count[31], temp_count[30], temp_count[29], temp_count[28], 
        temp_count[27], temp_count[26], temp_count[25], temp_count[24], 
        temp_count[23], temp_count[22], temp_count[21], temp_count[20], 
        temp_count[19], temp_count[18], temp_count[17], temp_count[16], 
        temp_count[15], temp_count[14], temp_count[13], temp_count[12], 
        temp_count[11], temp_count[10], temp_count[9], temp_count[8], 
        temp_count[7], temp_count[6], temp_count[5], temp_count[4], 
        temp_count[3], temp_count[2], temp_count[1], temp_count[0]}), 
        .dds_sin({dds_sin[7], dds_sin[6], dds_sin[5], dds_sin[4], 
        dds_sin[3], dds_sin[2], dds_sin[1], dds_sin[0]}), .dds_cos({
        dds_cos[7], dds_cos[6], dds_cos[5], dds_cos[4], dds_cos[3], 
        dds_cos[2], dds_cos[1], dds_cos[0]}), .IICE_comm2iice({
        \IICE_comm2iice[11] , \IICE_comm2iice[10] , 
        \IICE_comm2iice[9] , \IICE_comm2iice[8] , \IICE_comm2iice[7] , 
        \IICE_comm2iice[6] , \IICE_comm2iice[5] , \IICE_comm2iice[4] , 
        \IICE_comm2iice[3] , \IICE_comm2iice[2] , \IICE_comm2iice[1] , 
        \IICE_comm2iice[0] }), .freq_2(freq_2), .freq_14(freq_14), 
        .freq_15(freq_15), .freq_0(freq_0), .freq_1(freq_1), .freq_6(
        freq_6), .freq_10(freq_10), .freq_11(freq_11), .freq_13(
        freq_13), .BW_clk_c(BW_clk_c), .clk_dac2(clk_dac2), 
        .dac1_clk_c(dac1_clk_c), .temp_sck_c(temp_sck_c), .temp1_csn_c(
        temp1_csn_c), .temp2_csn_c(temp2_csn_c), .temp3_csn_c(
        temp3_csn_c), .temp_so_c(temp_so_c), .IICE_iice2comm(
        IICE_iice2comm));
    GND GND (.Y(GND_net_1));
    comm_block_x comm_block_INST (.IICE_comm2iice({\IICE_comm2iice[0] , 
        \IICE_comm2iice[1] , \IICE_comm2iice[2] , \IICE_comm2iice[3] , 
        \IICE_comm2iice[4] , \IICE_comm2iice[5] , \IICE_comm2iice[6] , 
        \IICE_comm2iice[7] , \IICE_comm2iice[8] , \IICE_comm2iice[9] , 
        \IICE_comm2iice[10] , \IICE_comm2iice[11] }), .IICE_iice2comm(
        IICE_iice2comm), .atck(atck), .atdi(atdi), .atdo(atdo), .atms(
        atms), .atrstb(atrstb));
    
endmodule


module build_sb_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module build_sb_CCC_0_FCCC(
       BW_clk_c,
       BW_clk_c_i_0,
       temp_sck_c,
       temp_sck_c_i_0,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output BW_clk_c;
output BW_clk_c_i_0;
output temp_sck_c;
output temp_sck_c_i_0;
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL2_net, GL1_net, VCC_net_1, GND_net_1;
    
    CLKINT GL1_INST (.A(GL1_net), .Y(temp_sck_c));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  GL1_INST_RNI8343 (.A(temp_sck_c), .Y(
        temp_sck_c_i_0));
    GND GND (.Y(GND_net_1));
    CLKINT GL2_INST (.A(GL2_net), .Y(BW_clk_c));
    CCC #( .INIT(210'h0000007FB8000044564003F0BC2B09C20E739DEFFC4C980C00B01)
        , .VCOFREQUENCY(600.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(), 
        .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(VCC_net_1), 
        .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), .NGMUX1_SEL(
        GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(GND_net_1), 
        .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(VCC_net_1), 
        .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(VCC_net_1), 
        .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(VCC_net_1), 
        .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(VCC_net_1), 
        .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(), .GL1(GL1_net), .GL2(
        GL2_net), .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    CFG1 #( .INIT(2'h1) )  GL2_INST_RNI98ED (.A(BW_clk_c), .Y(
        BW_clk_c_i_0));
    
endmodule


module build_sb(
       BW_clk_c,
       BW_clk_c_i_0,
       temp_sck_c,
       temp_sck_c_i_0
    );
output BW_clk_c;
output BW_clk_c_i_0;
output temp_sck_c;
output temp_sck_c_i_0;

    wire FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, GND_net_1, 
        VCC_net_1;
    
    build_sb_FABOSC_0_OSC FABOSC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    build_sb_CCC_0_FCCC CCC_0 (.BW_clk_c(BW_clk_c), .BW_clk_c_i_0(
        BW_clk_c_i_0), .temp_sck_c(temp_sck_c), .temp_sck_c_i_0(
        temp_sck_c_i_0), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    GND GND (.Y(GND_net_1));
    
endmodule


module build(
       BW,
       SENSE_DIN,
       adc_d0,
       BW_out,
       SENSE_DOUT,
       dac1_db,
       fl_a,
       fl_dq,
       ANTF_n1,
       ANTF_n2,
       DEVRST_N,
       GPIO10,
       GPIO11,
       GPIO8,
       GPIO9,
       GPS1_I0,
       GPS1_I1,
       GPS1_LD,
       GPS1_Q0,
       GPS1_Q1,
       GPS2_LD,
       GPS2_Q0,
       GPS2_Q1,
       GPS_I0,
       GPS_I1,
       adc_clk,
       adc_oen,
       adc_of,
       osc_vcc,
       temp_so,
       AMP_EN,
       BW_36,
       BW_clk,
       CSN_n1,
       CTR1,
       CTR2,
       CTR3,
       CTR4,
       CTR5,
       CTR6,
       CTR7,
       GPIO1,
       GPIO12,
       GPIO14,
       GPIO15,
       GPIO16,
       GPIO17,
       GPIO19,
       GPIO2,
       GPIO20,
       GPIO3,
       GPIO4,
       GPIO5,
       GPIO6,
       GPIO7,
       GPS1_IDLE,
       GPS1_PGM,
       GPS1_SCLK,
       GPS1_SDATA,
       GPS1_SHDN,
       REF_CE,
       REF_CLK,
       REF_DATA,
       REF_LD,
       REF_LE,
       REF_MXOUT,
       SENSE_CS_1,
       adc_shdn,
       clk_out_n1,
       clk_out_n2,
       dac1_clk,
       dac1_sleep,
       dac2_clk,
       dsa_clk,
       dsa_data,
       dsa_le,
       en_modul,
       fl_byten,
       fl_cen,
       fl_oen,
       fl_resetn,
       fl_ryby,
       fl_wen,
       fl_wpn,
       oclk_1,
       out1,
       out2,
       sr_cs1n,
       sr_cs2,
       sr_lbn,
       sr_oen,
       sr_ubn,
       sr_wen,
       temp1_csn,
       temp2_csn,
       temp3_csn,
       temp_sck,
       atck,
       atdi,
       atdo,
       atms,
       atrstb
    );
input  [14:0] BW;
input  [1:0] SENSE_DIN;
input  [13:0] adc_d0;
output [14:0] BW_out;
output [1:0] SENSE_DOUT;
output [13:5] dac1_db;
output [25:0] fl_a;
output [7:0] fl_dq;
input  ANTF_n1;
input  ANTF_n2;
input  DEVRST_N;
input  GPIO10;
input  GPIO11;
input  GPIO8;
input  GPIO9;
input  GPS1_I0;
input  GPS1_I1;
input  GPS1_LD;
input  GPS1_Q0;
input  GPS1_Q1;
input  GPS2_LD;
input  GPS2_Q0;
input  GPS2_Q1;
input  GPS_I0;
input  GPS_I1;
input  adc_clk;
input  adc_oen;
input  adc_of;
input  osc_vcc;
input  temp_so;
output AMP_EN;
output BW_36;
output BW_clk;
output CSN_n1;
output CTR1;
output CTR2;
output CTR3;
output CTR4;
output CTR5;
output CTR6;
output CTR7;
output GPIO1;
output GPIO12;
output GPIO14;
output GPIO15;
output GPIO16;
output GPIO17;
output GPIO19;
output GPIO2;
output GPIO20;
output GPIO3;
output GPIO4;
output GPIO5;
output GPIO6;
output GPIO7;
output GPS1_IDLE;
output GPS1_PGM;
output GPS1_SCLK;
output GPS1_SDATA;
output GPS1_SHDN;
output REF_CE;
output REF_CLK;
output REF_DATA;
output REF_LD;
output REF_LE;
output REF_MXOUT;
output SENSE_CS_1;
output adc_shdn;
output clk_out_n1;
output clk_out_n2;
output dac1_clk;
output dac1_sleep;
output dac2_clk;
output dsa_clk;
output dsa_data;
output dsa_le;
output en_modul;
output fl_byten;
output fl_cen;
output fl_oen;
output fl_resetn;
output fl_ryby;
output fl_wen;
output fl_wpn;
output oclk_1;
output out1;
output out2;
output sr_cs1n;
output sr_cs2;
output sr_lbn;
output sr_oen;
output sr_ubn;
output sr_wen;
output temp1_csn;
output temp2_csn;
output temp3_csn;
output temp_sck;
input  atck;
input  atdi;
output atdo;
input  atms;
input  atrstb;

    wire VCC_net_1, GND_net_1, \freq[7] , \freq[8] , \freq[9] , 
        \freq[13] , \freq[17] , \freq[18] , \freq[20] , \freq[21] , 
        \freq[22] , \temp_count_data[0] , \temp_count_data[1] , 
        \temp_count_data[2] , \temp_count_data[3] , 
        \temp_count_data[4] , \temp_count[0] , \temp_count[1] , 
        \temp_count[2] , \temp_count[3] , \temp_count[4] , 
        \temp_count[5] , \temp_count[6] , \temp_count[7] , 
        \temp_count[8] , \temp_count[9] , \temp_count[10] , 
        \temp_count[11] , \temp_count[12] , \temp_count[13] , 
        \temp_count[14] , \temp_count[15] , \temp_count[16] , 
        \temp_count[17] , \temp_count[18] , \temp_count[20] , 
        \temp_count[21] , \temp_count[22] , \temp_count[23] , 
        \temp_count[24] , \temp_count[25] , \temp_count[26] , 
        \temp_count[27] , \temp_count[28] , \temp_count[29] , 
        \temp_count[30] , \temp_count[31] , \temp3[0] , \temp3[1] , 
        \temp3[2] , \temp3[3] , \temp3[4] , \temp3[5] , \temp3[6] , 
        \temp3[7] , \temp3[8] , \temp3[9] , \temp3[10] , \temp3[11] , 
        \temp3[12] , \temp3[13] , \temp3[14] , \temp3[15] , \temp2[0] , 
        \temp2[1] , \temp2[2] , \temp2[3] , \temp2[4] , \temp2[5] , 
        \temp2[6] , \temp2[7] , \temp2[8] , \temp2[9] , \temp2[10] , 
        \temp2[11] , \temp2[12] , \temp2[13] , \temp2[14] , 
        \temp2[15] , \temp1[0] , \temp1[1] , \temp1[2] , \temp1[3] , 
        \temp1[4] , \temp1[5] , \temp1[6] , \temp1[7] , \temp1[8] , 
        \temp1[9] , \temp1[10] , \temp1[11] , \temp1[12] , \temp1[13] , 
        \temp1[14] , \temp1[15] , \sdv_count[0] , \sdv_count[1] , 
        \fr_adc_count[1] , \fr_adc_count[2] , \fr_adc_count[3] , 
        \fpga_shift_2[0] , \fpga_shift_2[1] , \fpga_shift_2[2] , 
        \fpga_shift_2[3] , \fpga_shift_2[4] , \fpga_shift_2[5] , 
        \fpga_shift_2[6] , \fpga_shift_2[7] , \fpga_shift_2[8] , 
        \fpga_shift_2[9] , \fpga_shift_2[10] , \fpga_shift_2[11] , 
        \fpga_shift_2[12] , \fpga_shift_2[13] , \fpga_shift_2[14] , 
        \fpga_count[0] , \dds_sin[0] , \dds_sin[1] , \dds_sin[2] , 
        \dds_sin[3] , \dds_sin[4] , \dds_sin[5] , \dds_sin[6] , 
        \dds_sin[7] , \dds_cos[0] , \dds_cos[1] , \dds_cos[2] , 
        \dds_cos[3] , \dds_cos[4] , \dds_cos[5] , \dds_cos[6] , 
        \dds_cos[7] , \data_from_adc[0][0] , \data_from_adc[0][1] , 
        \data_from_adc[0][2] , \data_from_adc[0][3] , 
        \data_from_adc[0][4] , \data_from_adc[0][5] , 
        \data_from_adc[0][6] , \data_from_adc[0][7] , 
        \data_from_adc[0][8] , \data_from_adc[0][9] , 
        \data_from_adc[0][10] , \data_from_adc[0][11] , 
        \data_from_adc[1][0] , \data_from_adc[1][1] , 
        \data_from_adc[1][2] , \data_from_adc[1][3] , 
        \data_from_adc[1][4] , \data_from_adc[1][5] , 
        \data_from_adc[1][6] , \data_from_adc[1][7] , 
        \data_from_adc[1][8] , \data_from_adc[1][9] , 
        \data_from_adc[1][10] , \data_from_adc[1][11] , 
        \data_from_adc[2][0] , \data_from_adc[2][1] , 
        \data_from_adc[2][2] , \data_from_adc[2][3] , 
        \data_from_adc[2][4] , \data_from_adc[2][5] , 
        \data_from_adc[2][6] , \data_from_adc[2][7] , 
        \data_from_adc[2][8] , \data_from_adc[2][9] , 
        \data_from_adc[2][10] , \data_from_adc[2][11] , 
        \data_from_adc[3][0] , \data_from_adc[3][1] , 
        \data_from_adc[3][2] , \data_from_adc[3][3] , 
        \data_from_adc[3][4] , \data_from_adc[3][5] , 
        \data_from_adc[3][6] , \data_from_adc[3][7] , 
        \data_from_adc[3][8] , \data_from_adc[3][9] , 
        \data_from_adc[3][10] , \data_from_adc[3][11] , 
        \data_from_adc[4][0] , \data_from_adc[4][1] , 
        \data_from_adc[4][2] , \data_from_adc[4][3] , 
        \data_from_adc[4][4] , \data_from_adc[4][5] , 
        \data_from_adc[4][6] , \data_from_adc[4][7] , 
        \data_from_adc[4][8] , \data_from_adc[4][9] , 
        \data_from_adc[4][10] , \data_from_adc[4][11] , 
        \data_from_adc[5][0] , \data_from_adc[5][1] , 
        \data_from_adc[5][2] , \data_from_adc[5][3] , 
        \data_from_adc[5][4] , \data_from_adc[5][5] , 
        \data_from_adc[5][6] , \data_from_adc[5][7] , 
        \data_from_adc[5][8] , \data_from_adc[5][9] , 
        \data_from_adc[5][10] , \data_from_adc[5][11] , 
        \data_from_adc[6][0] , \data_from_adc[6][1] , 
        \data_from_adc[6][2] , \data_from_adc[6][3] , 
        \data_from_adc[6][4] , \data_from_adc[6][5] , 
        \data_from_adc[6][6] , \data_from_adc[6][7] , 
        \data_from_adc[6][8] , \data_from_adc[6][9] , 
        \data_from_adc[6][10] , \data_from_adc[6][11] , 
        \data_from_adc[7][0] , \data_from_adc[7][1] , 
        \data_from_adc[7][2] , \data_from_adc[7][3] , 
        \data_from_adc[7][4] , \data_from_adc[7][5] , 
        \data_from_adc[7][6] , \data_from_adc[7][7] , 
        \data_from_adc[7][8] , \data_from_adc[7][9] , 
        \data_from_adc[7][10] , \data_from_adc[7][11] , 
        \data_from_adc[8][0] , \data_from_adc[8][1] , 
        \data_from_adc[8][2] , \data_from_adc[8][3] , 
        \data_from_adc[8][4] , \data_from_adc[8][5] , 
        \data_from_adc[8][6] , \data_from_adc[8][7] , 
        \data_from_adc[8][8] , \data_from_adc[8][9] , 
        \data_from_adc[8][10] , \data_from_adc[8][11] , \dac_count[1] , 
        \dac_count[2] , \dac_count[3] , \dac_count[4] , \dac_count[5] , 
        clk_dac2, ANTF_n1_c, ANTF_n2_c, \BW_c[0] , \BW_c[1] , 
        \BW_c[2] , \BW_c[3] , \BW_c[4] , \BW_c[5] , \BW_c[6] , 
        \BW_c[7] , \BW_c[8] , \BW_c[9] , \BW_c[10] , \BW_c[11] , 
        \BW_c[12] , \BW_c[13] , \BW_c[14] , GPIO10_c, GPIO11_c, 
        GPIO8_c, GPIO9_c, GPS1_I0_c, GPS1_I1_c, GPS1_LD_c, GPS1_Q0_c, 
        GPS1_Q1_c, GPS2_LD_c, GPS2_Q0_c, GPS2_Q1_c, GPS_I0_c, GPS_I1_c, 
        GPIO6_c, GPIO4_c, adc_clk_c, \adc_d0_c[0] , \adc_d0_c[1] , 
        \adc_d0_c[2] , \adc_d0_c[3] , \adc_d0_c[4] , \adc_d0_c[5] , 
        \adc_d0_c[6] , \adc_d0_c[7] , \adc_d0_c[8] , \adc_d0_c[9] , 
        \adc_d0_c[10] , \adc_d0_c[11] , \adc_d0_c[12] , \adc_d0_c[13] , 
        adc_oen_c, adc_of_c, osc_vcc_c, temp_so_c, BW_clk_c, 
        \BW_out_c[0] , \BW_out_c[1] , \BW_out_c[2] , \BW_out_c[3] , 
        \BW_out_c[4] , \BW_out_c[5] , \BW_out_c[6] , \BW_out_c[7] , 
        \BW_out_c[8] , \BW_out_c[9] , \BW_out_c[10] , \BW_out_c[11] , 
        \BW_out_c[12] , \BW_out_c[13] , \BW_out_c[14] , GPIO14_c, 
        GPIO16_c, GPIO3_c, GPIO5_c, GPIO7_c, SENSE_CS_1_c, 
        \SENSE_DOUT_c[1] , dac1_clk_c, \dac1_db_c[5] , \dac1_db_c[6] , 
        \dac1_db_c[7] , \dac1_db_c[8] , \dac1_db_c[9] , 
        \dac1_db_c[10] , \dac1_db_c[11] , \dac1_db_c[12] , 
        \dac1_db_c[13] , dac2_clk_c, oclk_1_c, temp1_csn_c, 
        temp2_csn_c, temp3_csn_c, temp_sck_c, \dac_count[6] , 
        \dac_count[7] , \fpga_count[1] , \fpga_count[2] , 
        \fpga_count[3] , \fpga_count[4] , \fpga_count[5] , 
        \fpga_count[6] , \fpga_count[7] , \fpga_count[8] , 
        \fpga_count[9] , \fpga_count[10] , \fpga_count[11] , 
        \fpga_count[12] , \fpga_count[13] , \fpga_count[14] , 
        BW_clk_c_i_0, temp_sck_c_i_0, GPIO9_c_i_0, GPIO8_c_i_0, 
        \temp_count[19] ;
    
    INBUF \BW_ibuf[9]  (.PAD(BW[9]), .Y(\BW_c[9] ));
    INBUF GPS1_I1_ibuf (.PAD(GPS1_I1), .Y(GPS1_I1_c));
    INBUF \BW_ibuf[3]  (.PAD(BW[3]), .Y(\BW_c[3] ));
    INBUF \adc_d0_ibuf[8]  (.PAD(adc_d0[8]), .Y(\adc_d0_c[8] ));
    TRIBUFF \fl_dq_obuft[1]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[1]));
    OUTBUF \BW_out_obuf[7]  (.D(\BW_out_c[7] ), .PAD(BW_out[7]));
    OUTBUF GPIO3_obuf (.D(GPIO3_c), .PAD(GPIO3));
    INBUF \adc_d0_ibuf[6]  (.PAD(adc_d0[6]), .Y(\adc_d0_c[6] ));
    INBUF \BW_ibuf[5]  (.PAD(BW[5]), .Y(\BW_c[5] ));
    OUTBUF \BW_out_obuf[8]  (.D(\BW_out_c[8] ), .PAD(BW_out[8]));
    INBUF GPS2_Q1_ibuf (.PAD(GPS2_Q1), .Y(GPS2_Q1_c));
    led_igloo led_igloo_0 (.sdv_count({\sdv_count[1] , \sdv_count[0] })
        , .temp_count_data({\temp_count_data[4] , \temp_count_data[3] , 
        \temp_count_data[2] , \temp_count_data[1] , 
        \temp_count_data[0] }), .BW_c({\BW_c[14] , \BW_c[13] , 
        \BW_c[12] , \BW_c[11] , \BW_c[10] , \BW_c[9] , \BW_c[8] , 
        \BW_c[7] , \BW_c[6] , \BW_c[5] , \BW_c[4] , \BW_c[3] , 
        \BW_c[2] , \BW_c[1] , \BW_c[0] }), .fpga_shift_2({
        \fpga_shift_2[14] , \fpga_shift_2[13] , \fpga_shift_2[12] , 
        \fpga_shift_2[11] , \fpga_shift_2[10] , \fpga_shift_2[9] , 
        \fpga_shift_2[8] , \fpga_shift_2[7] , \fpga_shift_2[6] , 
        \fpga_shift_2[5] , \fpga_shift_2[4] , \fpga_shift_2[3] , 
        \fpga_shift_2[2] , \fpga_shift_2[1] , \fpga_shift_2[0] }), 
        .BW_out_c({\BW_out_c[14] , \BW_out_c[13] , \BW_out_c[12] , 
        \BW_out_c[11] , \BW_out_c[10] , \BW_out_c[9] , \BW_out_c[8] , 
        \BW_out_c[7] , \BW_out_c[6] , \BW_out_c[5] , \BW_out_c[4] , 
        \BW_out_c[3] , \BW_out_c[2] , \BW_out_c[1] , \BW_out_c[0] }), 
        .fpga_count({\fpga_count[14] , \fpga_count[13] , 
        \fpga_count[12] , \fpga_count[11] , \fpga_count[10] , 
        \fpga_count[9] , \fpga_count[8] , \fpga_count[7] , 
        \fpga_count[6] , \fpga_count[5] , \fpga_count[4] , 
        \fpga_count[3] , \fpga_count[2] , \fpga_count[1] , 
        \fpga_count[0] }), .\data_from_adc[6] ({\data_from_adc[6][11] , 
        \data_from_adc[6][10] , \data_from_adc[6][9] , 
        \data_from_adc[6][8] , \data_from_adc[6][7] , 
        \data_from_adc[6][6] , \data_from_adc[6][5] , 
        \data_from_adc[6][4] , \data_from_adc[6][3] , 
        \data_from_adc[6][2] , \data_from_adc[6][1] , 
        \data_from_adc[6][0] }), .\data_from_adc[7] ({
        \data_from_adc[7][11] , \data_from_adc[7][10] , 
        \data_from_adc[7][9] , \data_from_adc[7][8] , 
        \data_from_adc[7][7] , \data_from_adc[7][6] , 
        \data_from_adc[7][5] , \data_from_adc[7][4] , 
        \data_from_adc[7][3] , \data_from_adc[7][2] , 
        \data_from_adc[7][1] , \data_from_adc[7][0] }), 
        .\data_from_adc[8] ({\data_from_adc[8][11] , 
        \data_from_adc[8][10] , \data_from_adc[8][9] , 
        \data_from_adc[8][8] , \data_from_adc[8][7] , 
        \data_from_adc[8][6] , \data_from_adc[8][5] , 
        \data_from_adc[8][4] , \data_from_adc[8][3] , 
        \data_from_adc[8][2] , \data_from_adc[8][1] , 
        \data_from_adc[8][0] }), .fr_adc_count({\fr_adc_count[3] , 
        \fr_adc_count[2] , \fr_adc_count[1] }), .temp3({\temp3[15] , 
        \temp3[14] , \temp3[13] , \temp3[12] , \temp3[11] , 
        \temp3[10] , \temp3[9] , \temp3[8] , \temp3[7] , \temp3[6] , 
        \temp3[5] , \temp3[4] , \temp3[3] , \temp3[2] , \temp3[1] , 
        \temp3[0] }), .dac1_db_c({\dac1_db_c[13] , \dac1_db_c[12] , 
        \dac1_db_c[11] , \dac1_db_c[10] , \dac1_db_c[9] , 
        \dac1_db_c[8] , \dac1_db_c[7] , \dac1_db_c[6] , \dac1_db_c[5] })
        , .\data_from_adc[0] ({\data_from_adc[0][11] , 
        \data_from_adc[0][10] , \data_from_adc[0][9] , 
        \data_from_adc[0][8] , \data_from_adc[0][7] , 
        \data_from_adc[0][6] , \data_from_adc[0][5] , 
        \data_from_adc[0][4] , \data_from_adc[0][3] , 
        \data_from_adc[0][2] , \data_from_adc[0][1] , 
        \data_from_adc[0][0] }), .\data_from_adc[1] ({
        \data_from_adc[1][11] , \data_from_adc[1][10] , 
        \data_from_adc[1][9] , \data_from_adc[1][8] , 
        \data_from_adc[1][7] , \data_from_adc[1][6] , 
        \data_from_adc[1][5] , \data_from_adc[1][4] , 
        \data_from_adc[1][3] , \data_from_adc[1][2] , 
        \data_from_adc[1][1] , \data_from_adc[1][0] }), 
        .\data_from_adc[3] ({\data_from_adc[3][11] , 
        \data_from_adc[3][10] , \data_from_adc[3][9] , 
        \data_from_adc[3][8] , \data_from_adc[3][7] , 
        \data_from_adc[3][6] , \data_from_adc[3][5] , 
        \data_from_adc[3][4] , \data_from_adc[3][3] , 
        \data_from_adc[3][2] , \data_from_adc[3][1] , 
        \data_from_adc[3][0] }), .\data_from_adc[2] ({
        \data_from_adc[2][11] , \data_from_adc[2][10] , 
        \data_from_adc[2][9] , \data_from_adc[2][8] , 
        \data_from_adc[2][7] , \data_from_adc[2][6] , 
        \data_from_adc[2][5] , \data_from_adc[2][4] , 
        \data_from_adc[2][3] , \data_from_adc[2][2] , 
        \data_from_adc[2][1] , \data_from_adc[2][0] }), 
        .\data_from_adc[4] ({\data_from_adc[4][11] , 
        \data_from_adc[4][10] , \data_from_adc[4][9] , 
        \data_from_adc[4][8] , \data_from_adc[4][7] , 
        \data_from_adc[4][6] , \data_from_adc[4][5] , 
        \data_from_adc[4][4] , \data_from_adc[4][3] , 
        \data_from_adc[4][2] , \data_from_adc[4][1] , 
        \data_from_adc[4][0] }), .\data_from_adc[5] ({
        \data_from_adc[5][11] , \data_from_adc[5][10] , 
        \data_from_adc[5][9] , \data_from_adc[5][8] , 
        \data_from_adc[5][7] , \data_from_adc[5][6] , 
        \data_from_adc[5][5] , \data_from_adc[5][4] , 
        \data_from_adc[5][3] , \data_from_adc[5][2] , 
        \data_from_adc[5][1] , \data_from_adc[5][0] }), .temp1({
        \temp1[15] , \temp1[14] , \temp1[13] , \temp1[12] , 
        \temp1[11] , \temp1[10] , \temp1[9] , \temp1[8] , \temp1[7] , 
        \temp1[6] , \temp1[5] , \temp1[4] , \temp1[3] , \temp1[2] , 
        \temp1[1] , \temp1[0] }), .temp2({\temp2[15] , \temp2[14] , 
        \temp2[13] , \temp2[12] , \temp2[11] , \temp2[10] , \temp2[9] , 
        \temp2[8] , \temp2[7] , \temp2[6] , \temp2[5] , \temp2[4] , 
        \temp2[3] , \temp2[2] , \temp2[1] , \temp2[0] }), 
        .SENSE_DOUT_c({\SENSE_DOUT_c[1] }), .dac_count({\dac_count[7] , 
        \dac_count[6] , \dac_count[5] , \dac_count[4] , \dac_count[3] , 
        \dac_count[2] , \dac_count[1] }), .temp_count({
        \temp_count[31] , \temp_count[30] , \temp_count[29] , 
        \temp_count[28] , \temp_count[27] , \temp_count[26] , 
        \temp_count[25] , \temp_count[24] , \temp_count[23] , 
        \temp_count[22] , \temp_count[21] , \temp_count[20] , 
        \temp_count[19] , \temp_count[18] , \temp_count[17] , 
        \temp_count[16] , \temp_count[15] , \temp_count[14] , 
        \temp_count[13] , \temp_count[12] , \temp_count[11] , 
        \temp_count[10] , \temp_count[9] , \temp_count[8] , 
        \temp_count[7] , \temp_count[6] , \temp_count[5] , 
        \temp_count[4] , \temp_count[3] , \temp_count[2] , 
        \temp_count[1] , \temp_count[0] }), .dds_cos({\dds_cos[7] , 
        \dds_cos[6] , \dds_cos[5] , \dds_cos[4] , \dds_cos[3] , 
        \dds_cos[2] , \dds_cos[1] , \dds_cos[0] }), .dds_sin({
        \dds_sin[7] , \dds_sin[6] , \dds_sin[5] , \dds_sin[4] , 
        \dds_sin[3] , \dds_sin[2] , \dds_sin[1] , \dds_sin[0] }), 
        .adc_d0_c({\adc_d0_c[13] , \adc_d0_c[12] , \adc_d0_c[11] , 
        \adc_d0_c[10] , \adc_d0_c[9] , \adc_d0_c[8] , \adc_d0_c[7] , 
        \adc_d0_c[6] , \adc_d0_c[5] , \adc_d0_c[4] , \adc_d0_c[3] , 
        \adc_d0_c[2] , \adc_d0_c[1] , \adc_d0_c[0] }), .freq_10(
        \freq[17] ), .freq_11(\freq[18] ), .freq_0(\freq[7] ), .freq_1(
        \freq[8] ), .freq_13(\freq[20] ), .freq_14(\freq[21] ), 
        .freq_15(\freq[22] ), .freq_6(\freq[13] ), .freq_2(\freq[9] ), 
        .temp_sck_c(temp_sck_c), .BW_clk_c_i_0(BW_clk_c_i_0), 
        .BW_clk_c(BW_clk_c), .GPIO4_c(GPIO4_c), .temp_sck_c_i_0(
        temp_sck_c_i_0), .temp_so_c(temp_so_c), .dac1_clk_c(dac1_clk_c)
        , .SENSE_CS_1_c(SENSE_CS_1_c), .GPIO16_c(GPIO16_c), .clk_dac2(
        clk_dac2), .GPIO14_c(GPIO14_c), .GPIO7_c(GPIO7_c), 
        .temp3_csn_c(temp3_csn_c), .temp2_csn_c(temp2_csn_c), 
        .temp1_csn_c(temp1_csn_c), .GPIO11_c(GPIO11_c), .oclk_1_c(
        oclk_1_c), .GPIO10_c(GPIO10_c), .dac2_clk_c(dac2_clk_c), 
        .adc_of_c(adc_of_c), .adc_oen_c(adc_oen_c), .adc_clk_c(
        adc_clk_c), .GPS_I1_c(GPS_I1_c), .GPS_I0_c(GPS_I0_c), 
        .GPS2_Q1_c(GPS2_Q1_c), .GPS2_Q0_c(GPS2_Q0_c), .GPS2_LD_c(
        GPS2_LD_c), .GPS1_Q1_c(GPS1_Q1_c), .GPS1_Q0_c(GPS1_Q0_c), 
        .GPS1_LD_c(GPS1_LD_c), .GPS1_I1_c(GPS1_I1_c), .GPS1_I0_c(
        GPS1_I0_c), .GPIO9_c(GPIO9_c), .GPIO6_c(GPIO6_c), .osc_vcc_c(
        osc_vcc_c), .ANTF_n2_c(ANTF_n2_c), .ANTF_n1_c(ANTF_n1_c), 
        .GPIO3_c(GPIO3_c), .GPIO5_c(GPIO5_c));
    TRIBUFF \fl_dq_obuft[7]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[7]));
    TRIBUFF \fl_dq_obuft[0]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[0]));
    OUTBUF \SENSE_DOUT_obuf[1]  (.D(\SENSE_DOUT_c[1] ), .PAD(
        SENSE_DOUT[1]));
    TRIBUFF sr_lbn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_lbn));
    TRIBUFF \fl_a_obuft[21]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[21]));
    INBUF ANTF_n1_ibuf (.PAD(ANTF_n1), .Y(ANTF_n1_c));
    INBUF \BW_ibuf[14]  (.PAD(BW[14]), .Y(\BW_c[14] ));
    OUTBUF adc_shdn_obuf (.D(VCC_net_1), .PAD(adc_shdn));
    TRIBUFF GPIO1_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(GPIO1));
    OUTBUF \dac1_db_obuf[9]  (.D(\dac1_db_c[9] ), .PAD(dac1_db[9]));
    OUTBUF \dac1_db_obuf[11]  (.D(\dac1_db_c[11] ), .PAD(dac1_db[11]));
    OUTBUF \dac1_db_obuf[6]  (.D(\dac1_db_c[6] ), .PAD(dac1_db[6]));
    TRIBUFF \fl_a_obuft[23]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[23]));
    OUTBUF CTR5_obuf (.D(GND_net_1), .PAD(CTR5));
    TRIBUFF \fl_dq_obuft[6]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[6]));
    TRIBUFF fl_cen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_cen));
    OUTBUF \dac1_db_obuf[10]  (.D(\dac1_db_c[10] ), .PAD(dac1_db[10]));
    INBUF \adc_d0_ibuf[13]  (.PAD(adc_d0[13]), .Y(\adc_d0_c[13] ));
    INBUF \BW_ibuf[2]  (.PAD(BW[2]), .Y(\BW_c[2] ));
    TRIBUFF REF_LE_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_LE));
    INBUF \BW_ibuf[11]  (.PAD(BW[11]), .Y(\BW_c[11] ));
    OUTBUF out1_obuf (.D(GND_net_1), .PAD(out1));
    OUTBUF CTR3_obuf (.D(GND_net_1), .PAD(CTR3));
    INBUF adc_oen_ibuf (.PAD(adc_oen), .Y(adc_oen_c));
    TRIBUFF REF_MXOUT_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        REF_MXOUT));
    INBUF \adc_d0_ibuf[9]  (.PAD(adc_d0[9]), .Y(\adc_d0_c[9] ));
    INBUF GPS1_I0_ibuf (.PAD(GPS1_I0), .Y(GPS1_I0_c));
    INBUF \adc_d0_ibuf[1]  (.PAD(adc_d0[1]), .Y(\adc_d0_c[1] ));
    TRIBUFF \fl_a_obuft[10]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[10]));
    OUTBUF CTR1_obuf (.D(GND_net_1), .PAD(CTR1));
    GND GND (.Y(GND_net_1));
    INBUF \SENSE_DIN_ibuf[0]  (.PAD(SENSE_DIN[0]), .Y(GPIO6_c));
    INBUF GPS2_Q0_ibuf (.PAD(GPS2_Q0), .Y(GPS2_Q0_c));
    OUTBUF \BW_out_obuf[11]  (.D(\BW_out_c[11] ), .PAD(BW_out[11]));
    OUTBUF \BW_out_obuf[6]  (.D(\BW_out_c[6] ), .PAD(BW_out[6]));
    OUTBUF \BW_out_obuf[1]  (.D(\BW_out_c[1] ), .PAD(BW_out[1]));
    OUTBUF GPIO12_obuf (.D(VCC_net_1), .PAD(GPIO12));
    OUTBUF GPIO15_obuf (.D(GND_net_1), .PAD(GPIO15));
    TRIBUFF \fl_a_obuft[17]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[17]));
    OUTBUF GPIO19_obuf (.D(GND_net_1), .PAD(GPIO19));
    TRIBUFF sr_cs2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_cs2));
    INBUF osc_vcc_ibuf (.PAD(osc_vcc), .Y(osc_vcc_c));
    syn_identify_core0_0 ident_coreinst (.BW_c({\BW_c[14] , \BW_c[13] , 
        \BW_c[12] , \BW_c[11] , \BW_c[10] , \BW_c[9] , \BW_c[8] , 
        \BW_c[7] , \BW_c[6] , \BW_c[5] , \BW_c[4] , \BW_c[3] , 
        \BW_c[2] , \BW_c[1] , \BW_c[0] }), .BW_out_c({\BW_out_c[14] , 
        \BW_out_c[13] , \BW_out_c[12] , \BW_out_c[11] , \BW_out_c[10] , 
        \BW_out_c[9] , \BW_out_c[8] , \BW_out_c[7] , \BW_out_c[6] , 
        \BW_out_c[5] , \BW_out_c[4] , \BW_out_c[3] , \BW_out_c[2] , 
        \BW_out_c[1] , \BW_out_c[0] }), .dac_count({\dac_count[7] , 
        \dac_count[6] , \dac_count[5] , \dac_count[4] , \dac_count[3] , 
        \dac_count[2] , \dac_count[1] }), .dac1_db_c({\dac1_db_c[13] , 
        \dac1_db_c[12] , \dac1_db_c[11] , \dac1_db_c[10] , 
        \dac1_db_c[9] , \dac1_db_c[8] , \dac1_db_c[7] , \dac1_db_c[6] , 
        \dac1_db_c[5] }), .\data_from_adc[8] ({\data_from_adc[8][11] , 
        \data_from_adc[8][10] , \data_from_adc[8][9] , 
        \data_from_adc[8][8] , \data_from_adc[8][7] , 
        \data_from_adc[8][6] , \data_from_adc[8][5] , 
        \data_from_adc[8][4] , \data_from_adc[8][3] , 
        \data_from_adc[8][2] , \data_from_adc[8][1] , 
        \data_from_adc[8][0] }), .\data_from_adc[7] ({
        \data_from_adc[7][11] , \data_from_adc[7][10] , 
        \data_from_adc[7][9] , \data_from_adc[7][8] , 
        \data_from_adc[7][7] , \data_from_adc[7][6] , 
        \data_from_adc[7][5] , \data_from_adc[7][4] , 
        \data_from_adc[7][3] , \data_from_adc[7][2] , 
        \data_from_adc[7][1] , \data_from_adc[7][0] }), 
        .\data_from_adc[6] ({\data_from_adc[6][11] , 
        \data_from_adc[6][10] , \data_from_adc[6][9] , 
        \data_from_adc[6][8] , \data_from_adc[6][7] , 
        \data_from_adc[6][6] , \data_from_adc[6][5] , 
        \data_from_adc[6][4] , \data_from_adc[6][3] , 
        \data_from_adc[6][2] , \data_from_adc[6][1] , 
        \data_from_adc[6][0] }), .\data_from_adc[4] ({
        \data_from_adc[4][11] , \data_from_adc[4][10] , 
        \data_from_adc[4][9] , \data_from_adc[4][8] , 
        \data_from_adc[4][7] , \data_from_adc[4][6] , 
        \data_from_adc[4][5] , \data_from_adc[4][4] , 
        \data_from_adc[4][3] , \data_from_adc[4][2] , 
        \data_from_adc[4][1] , \data_from_adc[4][0] }), 
        .\data_from_adc[5] ({\data_from_adc[5][11] , 
        \data_from_adc[5][10] , \data_from_adc[5][9] , 
        \data_from_adc[5][8] , \data_from_adc[5][7] , 
        \data_from_adc[5][6] , \data_from_adc[5][5] , 
        \data_from_adc[5][4] , \data_from_adc[5][3] , 
        \data_from_adc[5][2] , \data_from_adc[5][1] , 
        \data_from_adc[5][0] }), .\data_from_adc[3] ({
        \data_from_adc[3][11] , \data_from_adc[3][10] , 
        \data_from_adc[3][9] , \data_from_adc[3][8] , 
        \data_from_adc[3][7] , \data_from_adc[3][6] , 
        \data_from_adc[3][5] , \data_from_adc[3][4] , 
        \data_from_adc[3][3] , \data_from_adc[3][2] , 
        \data_from_adc[3][1] , \data_from_adc[3][0] }), 
        .\data_from_adc[2] ({\data_from_adc[2][11] , 
        \data_from_adc[2][10] , \data_from_adc[2][9] , 
        \data_from_adc[2][8] , \data_from_adc[2][7] , 
        \data_from_adc[2][6] , \data_from_adc[2][5] , 
        \data_from_adc[2][4] , \data_from_adc[2][3] , 
        \data_from_adc[2][2] , \data_from_adc[2][1] , 
        \data_from_adc[2][0] }), .\data_from_adc[1] ({
        \data_from_adc[1][11] , \data_from_adc[1][10] , 
        \data_from_adc[1][9] , \data_from_adc[1][8] , 
        \data_from_adc[1][7] , \data_from_adc[1][6] , 
        \data_from_adc[1][5] , \data_from_adc[1][4] , 
        \data_from_adc[1][3] , \data_from_adc[1][2] , 
        \data_from_adc[1][1] , \data_from_adc[1][0] }), 
        .\data_from_adc[0] ({\data_from_adc[0][11] , 
        \data_from_adc[0][10] , \data_from_adc[0][9] , 
        \data_from_adc[0][8] , \data_from_adc[0][7] , 
        \data_from_adc[0][6] , \data_from_adc[0][5] , 
        \data_from_adc[0][4] , \data_from_adc[0][3] , 
        \data_from_adc[0][2] , \data_from_adc[0][1] , 
        \data_from_adc[0][0] }), .fpga_count({\fpga_count[14] , 
        \fpga_count[13] , \fpga_count[12] , \fpga_count[11] , 
        \fpga_count[10] , \fpga_count[9] , \fpga_count[8] , 
        \fpga_count[7] , \fpga_count[6] , \fpga_count[5] , 
        \fpga_count[4] , \fpga_count[3] , \fpga_count[2] , 
        \fpga_count[1] , \fpga_count[0] }), .fr_adc_count({
        \fr_adc_count[3] , \fr_adc_count[2] , \fr_adc_count[1] }), 
        .fpga_shift_2({\fpga_shift_2[14] , \fpga_shift_2[13] , 
        \fpga_shift_2[12] , \fpga_shift_2[11] , \fpga_shift_2[10] , 
        \fpga_shift_2[9] , \fpga_shift_2[8] , \fpga_shift_2[7] , 
        \fpga_shift_2[6] , \fpga_shift_2[5] , \fpga_shift_2[4] , 
        \fpga_shift_2[3] , \fpga_shift_2[2] , \fpga_shift_2[1] , 
        \fpga_shift_2[0] }), .sdv_count({\sdv_count[1] , 
        \sdv_count[0] }), .temp1({\temp1[15] , \temp1[14] , 
        \temp1[13] , \temp1[12] , \temp1[11] , \temp1[10] , \temp1[9] , 
        \temp1[8] , \temp1[7] , \temp1[6] , \temp1[5] , \temp1[4] , 
        \temp1[3] , \temp1[2] , \temp1[1] , \temp1[0] }), .temp2({
        \temp2[15] , \temp2[14] , \temp2[13] , \temp2[12] , 
        \temp2[11] , \temp2[10] , \temp2[9] , \temp2[8] , \temp2[7] , 
        \temp2[6] , \temp2[5] , \temp2[4] , \temp2[3] , \temp2[2] , 
        \temp2[1] , \temp2[0] }), .temp3({\temp3[15] , \temp3[14] , 
        \temp3[13] , \temp3[12] , \temp3[11] , \temp3[10] , \temp3[9] , 
        \temp3[8] , \temp3[7] , \temp3[6] , \temp3[5] , \temp3[4] , 
        \temp3[3] , \temp3[2] , \temp3[1] , \temp3[0] }), 
        .temp_count_data({\temp_count_data[4] , \temp_count_data[3] , 
        \temp_count_data[2] , \temp_count_data[1] , 
        \temp_count_data[0] }), .temp_count({\temp_count[31] , 
        \temp_count[30] , \temp_count[29] , \temp_count[28] , 
        \temp_count[27] , \temp_count[26] , \temp_count[25] , 
        \temp_count[24] , \temp_count[23] , \temp_count[22] , 
        \temp_count[21] , \temp_count[20] , \temp_count[19] , 
        \temp_count[18] , \temp_count[17] , \temp_count[16] , 
        \temp_count[15] , \temp_count[14] , \temp_count[13] , 
        \temp_count[12] , \temp_count[11] , \temp_count[10] , 
        \temp_count[9] , \temp_count[8] , \temp_count[7] , 
        \temp_count[6] , \temp_count[5] , \temp_count[4] , 
        \temp_count[3] , \temp_count[2] , \temp_count[1] , 
        \temp_count[0] }), .dds_sin({\dds_sin[7] , \dds_sin[6] , 
        \dds_sin[5] , \dds_sin[4] , \dds_sin[3] , \dds_sin[2] , 
        \dds_sin[1] , \dds_sin[0] }), .dds_cos({\dds_cos[7] , 
        \dds_cos[6] , \dds_cos[5] , \dds_cos[4] , \dds_cos[3] , 
        \dds_cos[2] , \dds_cos[1] , \dds_cos[0] }), .freq_2(\freq[9] ), 
        .freq_14(\freq[21] ), .freq_15(\freq[22] ), .freq_0(\freq[7] ), 
        .freq_1(\freq[8] ), .freq_6(\freq[13] ), .freq_10(\freq[17] ), 
        .freq_11(\freq[18] ), .freq_13(\freq[20] ), .atck(atck), .atdi(
        atdi), .atdo(atdo), .atms(atms), .atrstb(atrstb), .BW_clk_c(
        BW_clk_c), .clk_dac2(clk_dac2), .dac1_clk_c(dac1_clk_c), 
        .temp_sck_c(temp_sck_c), .temp1_csn_c(temp1_csn_c), 
        .temp2_csn_c(temp2_csn_c), .temp3_csn_c(temp3_csn_c), 
        .temp_so_c(temp_so_c));
    TRIBUFF dsa_le_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(dsa_le));
    INBUF \BW_ibuf[0]  (.PAD(BW[0]), .Y(\BW_c[0] ));
    TRIBUFF GPS1_SCLK_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_SCLK));
    TRIBUFF GPS1_PGM_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_PGM));
    TRIBUFF \fl_dq_obuft[3]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[3]));
    TRIBUFF \fl_a_obuft[12]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[12]));
    TRIBUFF GPS1_SHDN_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_SHDN));
    OUTBUF GPIO14_obuf (.D(GPIO14_c), .PAD(GPIO14));
    OUTBUF AMP_EN_obuf (.D(GND_net_1), .PAD(AMP_EN));
    INBUF \adc_d0_ibuf[3]  (.PAD(adc_d0[3]), .Y(\adc_d0_c[3] ));
    TRIBUFF \fl_a_obuft[15]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[15]));
    INBUF GPS1_Q1_ibuf (.PAD(GPS1_Q1), .Y(GPS1_Q1_c));
    OUTBUF \BW_out_obuf[10]  (.D(\BW_out_c[10] ), .PAD(BW_out[10]));
    TRIBUFF \SENSE_DOUT_obuft[0]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        SENSE_DOUT[0]));
    OUTBUF \BW_out_obuf[9]  (.D(\BW_out_c[9] ), .PAD(BW_out[9]));
    OUTBUF CTR4_obuf (.D(GND_net_1), .PAD(CTR4));
    VCC VCC (.Y(VCC_net_1));
    TRIBUFF fl_byten_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_byten));
    TRIBUFF \fl_a_obuft[0]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[0]));
    INBUF adc_clk_ibuf (.PAD(adc_clk), .Y(adc_clk_c));
    OUTBUF CTR2_obuf (.D(GND_net_1), .PAD(CTR2));
    TRIBUFF sr_ubn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_ubn));
    TRIBUFF dac1_sleep_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        dac1_sleep));
    TRIBUFF \fl_a_obuft[8]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[8]));
    TRIBUFF REF_CLK_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_CLK));
    TRIBUFF GPS1_IDLE_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_IDLE));
    TRIBUFF dsa_data_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        dsa_data));
    TRIBUFF en_modul_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        en_modul));
    INBUF \adc_d0_ibuf[11]  (.PAD(adc_d0[11]), .Y(\adc_d0_c[11] ));
    OUTBUF temp3_csn_obuf (.D(temp3_csn_c), .PAD(temp3_csn));
    TRIBUFF REF_DATA_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        REF_DATA));
    OUTBUF \dac1_db_obuf[8]  (.D(\dac1_db_c[8] ), .PAD(dac1_db[8]));
    TRIBUFF fl_oen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_oen));
    INBUF GPS1_LD_ibuf (.PAD(GPS1_LD), .Y(GPS1_LD_c));
    OUTBUF \dac1_db_obuf[5]  (.D(\dac1_db_c[5] ), .PAD(dac1_db[5]));
    INBUF \adc_d0_ibuf[10]  (.PAD(adc_d0[10]), .Y(\adc_d0_c[10] ));
    TRIBUFF \fl_a_obuft[20]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[20]));
    TRIBUFF CSN_n1_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(CSN_n1));
    INBUF GPS_I0_ibuf (.PAD(GPS_I0), .Y(GPS_I0_c));
    OUTBUF \BW_out_obuf[13]  (.D(\BW_out_c[13] ), .PAD(BW_out[13]));
    TRIBUFF \fl_a_obuft[4]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[4]));
    INBUF \adc_d0_ibuf[2]  (.PAD(adc_d0[2]), .Y(\adc_d0_c[2] ));
    OUTBUF CTR6_obuf (.D(GPIO8_c_i_0), .PAD(CTR6));
    INBUF GPS1_Q0_ibuf (.PAD(GPS1_Q0), .Y(GPS1_Q0_c));
    INBUF \BW_ibuf[6]  (.PAD(BW[6]), .Y(\BW_c[6] ));
    TRIBUFF \fl_dq_obuft[5]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[5]));
    CFG1 #( .INIT(2'h1) )  CTR7_obuf_RNO (.A(GPIO9_c), .Y(GPIO9_c_i_0));
    INBUF GPS2_LD_ibuf (.PAD(GPS2_LD), .Y(GPS2_LD_c));
    INBUF \BW_ibuf[10]  (.PAD(BW[10]), .Y(\BW_c[10] ));
    TRIBUFF fl_resetn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_resetn));
    OUTBUF \BW_out_obuf[12]  (.D(\BW_out_c[12] ), .PAD(BW_out[12]));
    OUTBUF GPIO6_obuf (.D(GPIO6_c), .PAD(GPIO6));
    TRIBUFF \fl_a_obuft[5]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[5]));
    TRIBUFF \fl_a_obuft[9]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[9]));
    CFG1 #( .INIT(2'h1) )  CTR6_obuf_RNO (.A(GPIO8_c), .Y(GPIO8_c_i_0));
    INBUF \BW_ibuf[8]  (.PAD(BW[8]), .Y(\BW_c[8] ));
    TRIBUFF fl_wen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_wen));
    TRIBUFF \fl_a_obuft[22]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[22]));
    TRIBUFF \fl_a_obuft[25]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[25]));
    OUTBUF BW_clk_obuf (.D(BW_clk_c), .PAD(BW_clk));
    TRIBUFF sr_oen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_oen));
    INBUF adc_of_ibuf (.PAD(adc_of), .Y(adc_of_c));
    INBUF GPIO9_ibuf (.PAD(GPIO9), .Y(GPIO9_c));
    INBUF GPIO8_ibuf (.PAD(GPIO8), .Y(GPIO8_c));
    TRIBUFF \fl_a_obuft[14]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[14]));
    TRIBUFF sr_wen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_wen));
    INBUF \adc_d0_ibuf[4]  (.PAD(adc_d0[4]), .Y(\adc_d0_c[4] ));
    OUTBUF GPIO20_obuf (.D(GND_net_1), .PAD(GPIO20));
    TRIBUFF BW_36_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(BW_36));
    TRIBUFF out2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(out2));
    OUTBUF \dac1_db_obuf[12]  (.D(\dac1_db_c[12] ), .PAD(dac1_db[12]));
    OUTBUF \BW_out_obuf[5]  (.D(\BW_out_c[5] ), .PAD(BW_out[5]));
    INBUF \BW_ibuf[12]  (.PAD(BW[12]), .Y(\BW_c[12] ));
    OUTBUF GPIO7_obuf (.D(GPIO7_c), .PAD(GPIO7));
    INBUF GPIO10_ibuf (.PAD(GPIO10), .Y(GPIO10_c));
    INBUF temp_so_ibuf (.PAD(temp_so), .Y(temp_so_c));
    TRIBUFF REF_CE_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_CE));
    INBUF \adc_d0_ibuf[0]  (.PAD(adc_d0[0]), .Y(\adc_d0_c[0] ));
    TRIBUFF \fl_a_obuft[18]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[18]));
    OUTBUF temp2_csn_obuf (.D(temp2_csn_c), .PAD(temp2_csn));
    OUTBUF CTR7_obuf (.D(GPIO9_c_i_0), .PAD(CTR7));
    TRIBUFF fl_wpn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_wpn));
    INBUF \adc_d0_ibuf[5]  (.PAD(adc_d0[5]), .Y(\adc_d0_c[5] ));
    TRIBUFF dsa_clk_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(dsa_clk));
    TRIBUFF GPS1_SDATA_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_SDATA));
    TRIBUFF \fl_dq_obuft[4]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[4]));
    OUTBUF \BW_out_obuf[14]  (.D(\BW_out_c[14] ), .PAD(BW_out[14]));
    OUTBUF \BW_out_obuf[0]  (.D(\BW_out_c[0] ), .PAD(BW_out[0]));
    TRIBUFF REF_LD_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_LD));
    TRIBUFF clk_out_n2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        clk_out_n2));
    INBUF ANTF_n2_ibuf (.PAD(ANTF_n2), .Y(ANTF_n2_c));
    OUTBUF GPIO16_obuf (.D(GPIO16_c), .PAD(GPIO16));
    OUTBUF GPIO5_obuf (.D(GPIO5_c), .PAD(GPIO5));
    TRIBUFF \fl_a_obuft[11]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[11]));
    TRIBUFF \fl_a_obuft[19]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[19]));
    INBUF GPS_I1_ibuf (.PAD(GPS_I1), .Y(GPS_I1_c));
    TRIBUFF GPIO2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(GPIO2));
    INBUF \SENSE_DIN_ibuf[1]  (.PAD(SENSE_DIN[1]), .Y(GPIO4_c));
    build_sb build_sb_0 (.BW_clk_c(BW_clk_c), .BW_clk_c_i_0(
        BW_clk_c_i_0), .temp_sck_c(temp_sck_c), .temp_sck_c_i_0(
        temp_sck_c_i_0));
    TRIBUFF \fl_a_obuft[6]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[6]));
    INBUF \BW_ibuf[7]  (.PAD(BW[7]), .Y(\BW_c[7] ));
    INBUF \adc_d0_ibuf[7]  (.PAD(adc_d0[7]), .Y(\adc_d0_c[7] ));
    TRIBUFF fl_ryby_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_ryby));
    TRIBUFF \fl_a_obuft[13]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[13]));
    OUTBUF \dac1_db_obuf[7]  (.D(\dac1_db_c[7] ), .PAD(dac1_db[7]));
    OUTBUF GPIO4_obuf (.D(GPIO4_c), .PAD(GPIO4));
    OUTBUF temp1_csn_obuf (.D(temp1_csn_c), .PAD(temp1_csn));
    TRIBUFF \fl_a_obuft[1]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[1]));
    TRIBUFF \fl_a_obuft[3]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[3]));
    OUTBUF \dac1_db_obuf[13]  (.D(\dac1_db_c[13] ), .PAD(dac1_db[13]));
    TRIBUFF \fl_a_obuft[24]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[24]));
    INBUF \BW_ibuf[4]  (.PAD(BW[4]), .Y(\BW_c[4] ));
    INBUF \BW_ibuf[1]  (.PAD(BW[1]), .Y(\BW_c[1] ));
    OUTBUF temp_sck_obuf (.D(temp_sck_c), .PAD(temp_sck));
    TRIBUFF clk_out_n1_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        clk_out_n1));
    TRIBUFF \fl_a_obuft[16]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[16]));
    TRIBUFF \fl_dq_obuft[2]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[2]));
    INBUF \BW_ibuf[13]  (.PAD(BW[13]), .Y(\BW_c[13] ));
    TRIBUFF \fl_a_obuft[7]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[7]));
    OUTBUF oclk_1_obuf (.D(oclk_1_c), .PAD(oclk_1));
    OUTBUF dac1_clk_obuf (.D(dac1_clk_c), .PAD(dac1_clk));
    OUTBUF \BW_out_obuf[2]  (.D(\BW_out_c[2] ), .PAD(BW_out[2]));
    TRIBUFF GPIO17_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(GPIO17));
    TRIBUFF sr_cs1n_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_cs1n));
    OUTBUF \BW_out_obuf[4]  (.D(\BW_out_c[4] ), .PAD(BW_out[4]));
    TRIBUFF \fl_a_obuft[2]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[2]));
    OUTBUF dac2_clk_obuf (.D(dac2_clk_c), .PAD(dac2_clk));
    OUTBUF SENSE_CS_1_obuf (.D(SENSE_CS_1_c), .PAD(SENSE_CS_1));
    INBUF GPIO11_ibuf (.PAD(GPIO11), .Y(GPIO11_c));
    INBUF \adc_d0_ibuf[12]  (.PAD(adc_d0[12]), .Y(\adc_d0_c[12] ));
    OUTBUF \BW_out_obuf[3]  (.D(\BW_out_c[3] ), .PAD(BW_out[3]));
    
endmodule
