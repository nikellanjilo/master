`timescale 1 ns/100 ps
// Version: v11.6 SP1 11.6.1.6


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module led_igloo(
       temp_count_data,
       BW_out_c,
       BW_c,
       dac1_db_c,
       temp1,
       temp2,
       temp3,
       SENSE_DOUT_c,
       temp_count,
       adc_d0_c,
       freq_11,
       freq_2,
       freq_13,
       freq_14,
       freq_15,
       freq_0,
       freq_1,
       freq_10,
       freq_6,
       GPIO20_c,
       temp_sck_c,
       BW_clk_c,
       BW_clk_c_i_0,
       temp_so_c,
       GPIO4_c,
       temp_sck_c_i_0,
       dac1_clk_c,
       SENSE_CS_1_c,
       GPIO16_c,
       GPIO14_c,
       GPIO7_c,
       temp3_csn_c,
       temp2_csn_c,
       temp1_csn_c,
       GPIO11_c,
       GPIO10_c,
       dac2_clk_c,
       oclk_1_c,
       osc_vcc_c,
       adc_of_c,
       adc_oen_c,
       adc_clk_c,
       GPIO6_c,
       ANTF_n2_c,
       ANTF_n1_c,
       GPS1_LD_c,
       GPS1_I1_c,
       GPS1_I0_c,
       GPIO9_c,
       GPS2_Q0_c,
       GPS2_LD_c,
       GPS1_Q1_c,
       GPS1_Q0_c,
       GPS_I1_c,
       GPS_I0_c,
       GPS2_Q1_c,
       GPIO3_c,
       GPIO5_c
    );
output [4:0] temp_count_data;
output [14:0] BW_out_c;
input  [14:0] BW_c;
output [13:5] dac1_db_c;
output [15:0] temp1;
output [15:0] temp2;
output [15:0] temp3;
output [1:1] SENSE_DOUT_c;
output [31:0] temp_count;
input  [13:0] adc_d0_c;
output freq_11;
output freq_2;
output freq_13;
output freq_14;
output freq_15;
output freq_0;
output freq_1;
output freq_10;
output freq_6;
output GPIO20_c;
input  temp_sck_c;
input  BW_clk_c;
input  BW_clk_c_i_0;
input  temp_so_c;
input  GPIO4_c;
input  temp_sck_c_i_0;
output dac1_clk_c;
output SENSE_CS_1_c;
output GPIO16_c;
output GPIO14_c;
output GPIO7_c;
output temp3_csn_c;
output temp2_csn_c;
output temp1_csn_c;
input  GPIO11_c;
input  GPIO10_c;
output dac2_clk_c;
output oclk_1_c;
input  osc_vcc_c;
input  adc_of_c;
input  adc_oen_c;
input  adc_clk_c;
input  GPIO6_c;
input  ANTF_n2_c;
input  ANTF_n1_c;
input  GPS1_LD_c;
input  GPS1_I1_c;
input  GPS1_I0_c;
input  GPIO9_c;
input  GPS2_Q0_c;
input  GPS2_LD_c;
input  GPS1_Q1_c;
input  GPS1_Q0_c;
input  GPS_I1_c;
input  GPS_I0_c;
input  GPS2_Q1_c;
output GPIO3_c;
output GPIO5_c;

    wire \fpga_count[0]_net_1 , \fpga_count_s[0] , \dac_count_s[0] , 
        \cnt_freq[0]_net_1 , \cnt_freq_s[0] , \temp_state[0]_net_1 , 
        \temp_state_i_0[0] , \sdv_count[1]_net_1 , \sdv_count_i_0[1] , 
        \sdv_count[0]_net_1 , \sdv_count_i_0[0] , cnt_frame_0_sqmuxa, 
        N_333_i, temp_state26, N_322_i, fpga_flag_net_1, fpga_flag_i, 
        VCC_net_1, N_8_i_0, N_17_i_0, GND_net_1, N_6_i_0, N_113, 
        N_15_i_0, N_10_i_0, \fpga_shift_2[12]_net_1 , 
        \fpga_shift_2[13]_net_1 , \fpga_shift_2[14]_net_1 , 
        \fpga_data_receive[12]_net_1 , \fpga_data_receive[13]_net_1 , 
        \fpga_data_receive[14]_net_1 , \fpga_shift_2[0]_net_1 , 
        \fpga_shift_2[1]_net_1 , \fpga_shift_2[2]_net_1 , 
        \fpga_shift_2[3]_net_1 , \fpga_shift_2[4]_net_1 , 
        \fpga_shift_2[5]_net_1 , \fpga_shift_2[6]_net_1 , 
        \fpga_shift_2[7]_net_1 , \fpga_shift_2[8]_net_1 , 
        \fpga_shift_2[9]_net_1 , \fpga_shift_2[10]_net_1 , 
        \fpga_shift_2[11]_net_1 , \fpga_count[12]_net_1 , 
        \fpga_count[13]_net_1 , \fpga_count[14]_net_1 , 
        \fpga_data_receive[0]_net_1 , \fpga_data_receive[1]_net_1 , 
        \fpga_data_receive[2]_net_1 , \fpga_data_receive[3]_net_1 , 
        \fpga_data_receive[4]_net_1 , \fpga_data_receive[5]_net_1 , 
        \fpga_data_receive[6]_net_1 , \fpga_data_receive[7]_net_1 , 
        \fpga_data_receive[8]_net_1 , \fpga_data_receive[9]_net_1 , 
        \fpga_data_receive[10]_net_1 , \fpga_data_receive[11]_net_1 , 
        \temp_state[2]_net_1 , \temp_state_7[2] , \sdv_count_1[1] , 
        \fpga_count[1]_net_1 , \fpga_count[2]_net_1 , 
        \fpga_count[3]_net_1 , \fpga_count[4]_net_1 , 
        \fpga_count[5]_net_1 , \fpga_count[6]_net_1 , 
        \fpga_count[7]_net_1 , \fpga_count[8]_net_1 , 
        \fpga_count[9]_net_1 , \fpga_count[10]_net_1 , 
        \fpga_count[11]_net_1 , temp1_23, temp1_24, temp1_25, temp1_26, 
        N_726_i, N_719_i, N_712_i, N_705_i, N_698_i, N_691_i, N_684_i, 
        N_677_i, N_670_i, N_22_i_0, \temp_state[1]_net_1 , N_11_i_0, 
        temp2_40, temp2_41, temp2_42, temp1_11, temp1_12, temp1_13, 
        temp1_14, temp1_15, temp1_16, temp1_17, temp1_18, temp1_19, 
        temp1_20, temp1_21, temp1_22, temp3_57, temp3_58, temp2_27, 
        temp2_28, temp2_29, temp2_30, temp2_31, temp2_32, temp2_33, 
        temp2_34, temp2_35, temp2_36, temp2_37, temp2_38, temp2_39, 
        \data_from_adc[2][11]_net_1 , \data_from_adc[2]_70 , temp3_43, 
        temp3_44, temp3_45, temp3_46, temp3_47, temp3_48, temp3_49, 
        temp3_50, temp3_51, temp3_52, temp3_53, temp3_54, temp3_55, 
        temp3_56, \un1_data_from_adc[2]_1 , N_575_i_0, 
        \un1_data_from_adc[2]_1_i_0 , \data_from_adc[2][0]_net_1 , 
        \data_from_adc[2]_59 , \data_from_adc[2][1]_net_1 , 
        \data_from_adc[2]_60 , \data_from_adc[2][2]_net_1 , 
        \data_from_adc[2]_61 , \data_from_adc[2][3]_net_1 , 
        \data_from_adc[2]_62 , \data_from_adc[2][4]_net_1 , 
        \data_from_adc[2]_63 , \data_from_adc[2][5]_net_1 , 
        \data_from_adc[2]_64 , \data_from_adc[2][6]_net_1 , 
        \data_from_adc[2]_65 , \data_from_adc[2][7]_net_1 , 
        \data_from_adc[2]_66 , \data_from_adc[2][8]_net_1 , 
        \data_from_adc[2]_67 , \data_from_adc[2][9]_net_1 , 
        \data_from_adc[2]_68 , \data_from_adc[2][10]_net_1 , 
        \data_from_adc[2]_69 , freq15_i_0_net_1, N_445_i_0, 
        \un1_data_from_adc[2]_i_0 , \state[0]_net_1 , N_449_i_0, 
        N_70_i_0, \state[1]_net_1 , N_23_i_0, freq9_net_1, freq3, 
        freq3_i_0, clk_dac1_2_net_1, N_19_i_0, N_39_i_0, N_21, state15, 
        N_12_i_0, freq15_net_1, clk_dac2_net_1, cnt_freq6, 
        \cnt_freq[1]_net_1 , \cnt_freq_s[1] , \cnt_freq[2]_net_1 , 
        \cnt_freq_s[2] , \cnt_freq[3]_net_1 , \cnt_freq_s[3] , 
        \cnt_freq[4]_net_1 , \cnt_freq_s[4] , \cnt_freq[5]_net_1 , 
        \cnt_freq_s[5] , \cnt_freq[6]_net_1 , \cnt_freq_s[6] , 
        \cnt_freq[7]_net_1 , \cnt_freq_s[7] , \cnt_freq[8]_net_1 , 
        \cnt_freq_s[8] , \cnt_freq[9]_net_1 , \cnt_freq_s[9] , 
        \cnt_freq[10]_net_1 , \cnt_freq_s[10] , \cnt_freq[11]_net_1 , 
        \cnt_freq_s[11] , \cnt_freq[12]_net_1 , \cnt_freq_s[12] , 
        \cnt_freq[13]_net_1 , \cnt_freq_s[13] , \cnt_freq[14]_net_1 , 
        \cnt_freq_s[14] , \cnt_freq[15]_net_1 , \cnt_freq_s[15] , 
        \cnt_freq[16]_net_1 , \cnt_freq_s[16] , \cnt_freq[17]_net_1 , 
        \cnt_freq_s[17] , \cnt_freq[18]_net_1 , \cnt_freq_s[18] , 
        \cnt_freq[19]_net_1 , \cnt_freq_s[19] , \cnt_freq[20]_net_1 , 
        \cnt_freq_s[20] , \cnt_freq[21]_net_1 , \cnt_freq_s[21] , 
        \cnt_freq[22]_net_1 , \cnt_freq_s[22] , \cnt_freq[23]_net_1 , 
        \cnt_freq_s[23] , \cnt_freq[24]_net_1 , \cnt_freq_s[24] , 
        \cnt_freq[25]_net_1 , \cnt_freq_s[25] , \cnt_freq[26]_net_1 , 
        \cnt_freq_s[26] , \cnt_freq[27]_net_1 , \cnt_freq_s[27] , 
        \cnt_freq[28]_net_1 , \cnt_freq_s[28] , \cnt_freq[29]_net_1 , 
        \cnt_freq_s[29] , \cnt_freq[30]_net_1 , \cnt_freq_s[30] , 
        \cnt_freq[31]_net_1 , \cnt_freq_s[31]_net_1 , \cnt_s[0] , cnte, 
        \cnt[1]_net_1 , \cnt_s[1] , \cnt[2]_net_1 , \cnt_s[2] , 
        \cnt[3]_net_1 , \cnt_s[3] , \cnt[4]_net_1 , \cnt_s[4] , 
        \cnt[5]_net_1 , \cnt_s[5]_net_1 , \temp_count_s[0] , 
        \temp_count_s[1] , \temp_count_s[2] , \temp_count_s[3] , 
        \temp_count_s[4] , \temp_count_s[5] , \temp_count_s[6] , 
        \temp_count_s[7] , \temp_count_s[8] , \temp_count_s[9] , 
        \temp_count_s[10] , \temp_count_s[11] , \temp_count_s[12] , 
        \temp_count_s[13] , \temp_count_s[14] , \temp_count_s[15] , 
        \temp_count_s[16] , \temp_count_s[17] , \temp_count_s[18] , 
        \temp_count_s[19] , \temp_count_s[20] , \temp_count_s[21] , 
        \temp_count_s[22] , \temp_count_s[23] , \temp_count_s[24] , 
        \temp_count_s[25] , \temp_count_s[26] , \temp_count_s[27] , 
        \temp_count_s[28] , \temp_count_s[29] , \temp_count_s[30] , 
        \temp_count_s[31] , clk_dac14_net_1, \dac_count[1]_net_1 , 
        \dac_count_s[1] , \dac_count[2]_net_1 , \dac_count_s[2] , 
        \dac_count[3]_net_1 , \dac_count_s[3] , \dac_count[4]_net_1 , 
        \dac_count_s[4] , \dac_count[5]_net_1 , \dac_count_s[5] , 
        \dac_count[6]_net_1 , \dac_count_s[6] , \dac_count[7]_net_1 , 
        \dac_count_s[7] , \dac_count[8]_net_1 , \dac_count_s[8]_net_1 , 
        \fpga_count_s[1] , \fpga_count_s[2] , \fpga_count_s[3] , 
        \fpga_count_s[4] , \fpga_count_s[5] , \fpga_count_s[6] , 
        \fpga_count_s[7] , \fpga_count_s[8] , \fpga_count_s[9] , 
        \fpga_count_s[10] , \fpga_count_s[11] , \fpga_count_s[12] , 
        \fpga_count_s[13] , \fpga_count_s[14]_net_1 , fpga_flags, 
        temp3_csn_RNO_net_1, un1_temp_state_7_or, temp2_csn_1_sqmuxa, 
        temp2_csn_RNO_net_1, un1_temp_state29_3_or, 
        temp1_csn_RNO_net_1, un1_temp_state_8_or, \cnt_frame[3]_net_1 , 
        \cnt_frame_RNO[3]_net_1 , \cnt_frame_0_0_a2_0_2[3]_net_1 , 
        \cnt_frame[0]_net_1 , cnt_frame_1, \cnt_frame[1]_net_1 , 
        cnt_frame_0, \cnt_frame[2]_net_1 , cnt_frame, cnt_cry_cy, 
        N_36_i_0, \cnt_cry[0]_net_1 , \cnt_cry[1]_net_1 , 
        \cnt_cry[2]_net_1 , \cnt_cry[3]_net_1 , \cnt_cry[4]_net_1 , 
        temp_count_lcry_cy, temp_count_net_1, 
        temp_count6_cry_31_RNIPJ5K1_Y, temp_count6, 
        \temp_count_cry[0] , \temp_count_cry[1] , \temp_count_cry[2] , 
        \temp_count_cry[3] , \temp_count_cry[4] , \temp_count_cry[5] , 
        \temp_count_cry[6] , \temp_count_cry[7] , \temp_count_cry[8] , 
        \temp_count_cry[9] , \temp_count_cry[10] , 
        \temp_count_cry[11] , \temp_count_cry[12] , 
        \temp_count_cry[13] , \temp_count_cry[14] , 
        \temp_count_cry[15] , \temp_count_cry[16] , 
        \temp_count_cry[17] , \temp_count_cry[18] , 
        \temp_count_cry[19] , \temp_count_cry[20] , 
        \temp_count_cry[21] , \temp_count_cry[22] , 
        \temp_count_cry[23] , \temp_count_cry[24] , 
        \temp_count_cry[25] , \temp_count_cry[26] , 
        \temp_count_cry[27] , \temp_count_cry[28] , 
        \temp_count_cry[29] , \temp_count_cry[30] , 
        cnt_freq6_cry_7_net_1, cnt_freq6_cry_8_net_1, 
        cnt_freq6_cry_9_net_1, cnt_freq6_cry_10_net_1, 
        cnt_freq6_cry_11_net_1, cnt_freq6_cry_12_net_1, 
        cnt_freq6_cry_13_net_1, cnt_freq6_cry_14_net_1, 
        cnt_freq6_cry_15_net_1, cnt_freq6_cry_16_net_1, 
        cnt_freq6_cry_17_net_1, cnt_freq6_cry_18_net_1, 
        cnt_freq6_cry_19_net_1, cnt_freq6_cry_20_net_1, 
        cnt_freq6_cry_21_net_1, cnt_freq6_cry_22_net_1, 
        cnt_freq6_cry_23_net_1, cnt_freq6_cry_24_net_1, 
        cnt_freq6_cry_25_net_1, cnt_freq6_cry_26_net_1, 
        cnt_freq6_cry_27_net_1, cnt_freq6_cry_28_net_1, 
        cnt_freq6_cry_29_net_1, cnt_freq6_cry_30_net_1, 
        temp_count6_cry_7_net_1, temp_count6_cry_8_net_1, 
        temp_count6_cry_9_net_1, temp_count6_cry_10_net_1, 
        temp_count6_cry_11_net_1, temp_count6_cry_12_net_1, 
        temp_count6_cry_13_net_1, temp_count6_cry_14_net_1, 
        temp_count6_cry_15_net_1, temp_count6_cry_16_net_1, 
        temp_count6_cry_17_net_1, temp_count6_cry_18_net_1, 
        temp_count6_cry_19_net_1, temp_count6_cry_20_net_1, 
        temp_count6_cry_21_net_1, temp_count6_cry_22_net_1, 
        temp_count6_cry_23_net_1, temp_count6_cry_24_net_1, 
        temp_count6_cry_25_net_1, temp_count6_cry_26_net_1, 
        temp_count6_cry_27_net_1, temp_count6_cry_28_net_1, 
        temp_count6_cry_29_net_1, temp_count6_cry_30_net_1, 
        \fpga_flag4_0_data_tmp[0] , \fpga_flag4_0_data_tmp[1] , 
        \fpga_flag4_0_data_tmp[2] , \fpga_flag4_0_data_tmp[3] , 
        \fpga_flag4_0_data_tmp[4] , \fpga_flag4_0_data_tmp[5] , 
        \fpga_flag4_0_data_tmp[6] , fpga_count_s_459_FCO, 
        \fpga_count_cry[1]_net_1 , \fpga_count_cry[2]_net_1 , 
        \fpga_count_cry[3]_net_1 , \fpga_count_cry[4]_net_1 , 
        \fpga_count_cry[5]_net_1 , \fpga_count_cry[6]_net_1 , 
        \fpga_count_cry[7]_net_1 , \fpga_count_cry[8]_net_1 , 
        \fpga_count_cry[9]_net_1 , \fpga_count_cry[10]_net_1 , 
        \fpga_count_cry[11]_net_1 , \fpga_count_cry[12]_net_1 , 
        \fpga_count_cry[13]_net_1 , dac_count_s_460_FCO, 
        \dac_count_cry[1]_net_1 , \dac_count_cry[2]_net_1 , 
        \dac_count_cry[3]_net_1 , \dac_count_cry[4]_net_1 , 
        \dac_count_cry[5]_net_1 , \dac_count_cry[6]_net_1 , 
        \dac_count_cry[7]_net_1 , cnt_freq_s_461_FCO, 
        \cnt_freq_cry[1]_net_1 , \cnt_freq_cry[2]_net_1 , 
        \cnt_freq_cry[3]_net_1 , \cnt_freq_cry[4]_net_1 , 
        \cnt_freq_cry[5]_net_1 , \cnt_freq_cry[6]_net_1 , 
        \cnt_freq_cry[7]_net_1 , \cnt_freq_cry[8]_net_1 , 
        \cnt_freq_cry[9]_net_1 , \cnt_freq_cry[10]_net_1 , 
        \cnt_freq_cry[11]_net_1 , \cnt_freq_cry[12]_net_1 , 
        \cnt_freq_cry[13]_net_1 , \cnt_freq_cry[14]_net_1 , 
        \cnt_freq_cry[15]_net_1 , \cnt_freq_cry[16]_net_1 , 
        \cnt_freq_cry[17]_net_1 , \cnt_freq_cry[18]_net_1 , 
        \cnt_freq_cry[19]_net_1 , \cnt_freq_cry[20]_net_1 , 
        \cnt_freq_cry[21]_net_1 , \cnt_freq_cry[22]_net_1 , 
        \cnt_freq_cry[23]_net_1 , \cnt_freq_cry[24]_net_1 , 
        \cnt_freq_cry[25]_net_1 , \cnt_freq_cry[26]_net_1 , 
        \cnt_freq_cry[27]_net_1 , \cnt_freq_cry[28]_net_1 , 
        \cnt_freq_cry[29]_net_1 , \cnt_freq_cry[30]_net_1 , 
        \data_from_adc[2]_66_0_0_a2_0_out , 
        \data_from_adc[2]_66_0_0_a2_0_0 , N_22_i_1, 
        \un1_data_from_adc[2]lt10 , \un1_data_from_adc[2]_1lt10 , 
        freq3lt11, \data_from_adc[2]_66_0_0_a2_0 , 
        \data_from_adc[2]_59_0_0_a2_0 , 
        \SENSE_DOUT_2_1_u_i_a2_0[1]_net_1 , GPIO3_6_net_1, 
        \data_from_adc[2]_68_0_0_a2_0_out , 
        \data_from_adc[2]_59_0_0_a2_0_0 , N_183, N_76, N_58, N_182, 
        freq3lt8, N_178, \data_from_adc[2]_63_0_0_a2_0 , 
        \un1_data_from_adc[2]_2lto11_i_a2_7_net_1 , 
        \un1_data_from_adc[2]_2lto11_i_a2_6_net_1 , 
        \un1_data_from_adc[2]_2lto11_i_a2_5_net_1 , 
        \SENSE_DOUT_2_1_u_i_a2_0_0[1]_net_1 , freq3lto8_1_net_1, 
        GPIO3_9_net_1, GPIO3_8_net_1, GPIO3_7_net_1, GPIO5_13_net_1, 
        GPIO5_12_net_1, GPIO5_11_net_1, GPIO5_10_net_1, N_54, N_99, 
        \data_from_adc[2]_70_0_0_a2_0 , \data_from_adc[2]_68_0_0_a2_0 , 
        \un1_data_from_adc[2]lto8_0_net_1 , N_181, N_44, N_180, 
        \un1_data_from_adc[2]lt5 , N_109, \data_from_adc[2]_61_1 , 
        N_179, m10_0_0, \data_from_adc[2]_64_0_0_a2_1 , 
        \data_from_adc[2]_65_0_0_a2_1 , GPIO5_14_net_1, N_86, N_43, 
        N_80, N_3563_tz, N_52, \SENSE_DOUT_2_1_u_i_1[1]_net_1 ;
    
    ARI1 #( .INIT(20'h4AA00) )  dac_count_s_460 (.A(VCC_net_1), .B(
        GPIO20_c), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), .S(), 
        .Y(), .FCO(dac_count_s_460_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[11]  (.A(VCC_net_1), .B(
        \cnt_freq[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[10]_net_1 ), .S(\cnt_freq_s[11] ), .Y(), .FCO(
        \cnt_freq_cry[11]_net_1 ));
    CFG4 #( .INIT(16'h0051) )  freq9 (.A(\data_from_adc[2][11]_net_1 ), 
        .B(\data_from_adc[2][10]_net_1 ), .C(
        \un1_data_from_adc[2]lt10 ), .D(freq3), .Y(freq9_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[25]  (.A(VCC_net_1), .B(
        \cnt_freq[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[24]_net_1 ), .S(\cnt_freq_s[25] ), .Y(), .FCO(
        \cnt_freq_cry[25]_net_1 ));
    SLE \state[0]  (.D(N_449_i_0), .CLK(temp_sck_c_i_0), .EN(N_70_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  fpga_count_s_459 (.A(VCC_net_1), .B(
        \fpga_count[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(fpga_count_s_459_FCO));
    CFG2 #( .INIT(4'h1) )  \data_from_adc[2]_RNO_0[7]  (.A(
        \cnt[2]_net_1 ), .B(\cnt[1]_net_1 ), .Y(
        \data_from_adc[2]_66_0_0_a2_0 ));
    SLE \data_from_adc[2][6]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_65 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][6]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  GPIO5 (.A(GPIO5_14_net_1), .B(
        GPIO5_13_net_1), .C(GPIO5_12_net_1), .D(GPIO5_11_net_1), .Y(
        GPIO5_c));
    SLE \freq[17]  (.D(freq3_i_0), .CLK(temp_sck_c), .EN(N_575_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(freq_10));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_15 (.A(freq_0), .B(
        temp_count[15]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_14_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_15_net_1));
    CFG4 #( .INIT(16'h0010) )  temp1_23_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_76), .Y(temp1_23));
    SLE \fpga_count[2]  (.D(\fpga_count_s[2] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[2]_net_1 ));
    SLE \cnt_freq[26]  (.D(\cnt_freq_s[26] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[26]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_21 (.A(freq_14), .B(
        temp_count[21]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_20_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_21_net_1));
    CFG4 #( .INIT(16'h0800) )  temp3_43_0_0_a2 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(N_180));
    SLE \temp2[0]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_27), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[0]));
    CFG3 #( .INIT(8'h7F) )  freq3lto8_1 (.A(
        \data_from_adc[2][6]_net_1 ), .B(\data_from_adc[2][5]_net_1 ), 
        .C(\data_from_adc[2][4]_net_1 ), .Y(freq3lto8_1_net_1));
    SLE \dac1_db[13]  (.D(N_670_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[13]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIILLC9[3]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[3]), .D(
        GND_net_1), .FCI(\temp_count_cry[2] ), .S(\temp_count_s[3] ), 
        .Y(), .FCO(\temp_count_cry[3] ));
    CFG4 #( .INIT(16'h1000) )  temp3_58_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_178), .Y(temp3_58));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI75ACT[13]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[13]), .D(GND_net_1), .FCI(\temp_count_cry[12] ), .S(
        \temp_count_s[13] ), .Y(), .FCO(\temp_count_cry[13] ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_28 (.A(VCC_net_1), .B(
        temp_count[28]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_27_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_28_net_1));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_10 (.A(freq_0), .B(
        temp_count[10]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_9_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_10_net_1));
    SLE \cnt[0]  (.D(\cnt_s[0] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(GPIO7_c));
    SLE \temp1[13]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_24), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[13]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_14 (.A(VCC_net_1), .B(
        \cnt_freq[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_13_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_14_net_1));
    ARI1 #( .INIT(20'h45500) )  \cnt_cry_cy[0]  (.A(VCC_net_1), .B(
        N_36_i_0), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), .S(), 
        .Y(), .FCO(cnt_cry_cy));
    CFG1 #( .INIT(2'h1) )  fpga_flag_RNO (.A(fpga_flag_net_1), .Y(
        fpga_flag_i));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_39 (.A(
        \fpga_shift_2[3]_net_1 ), .B(\fpga_data_receive[2]_net_1 ), .C(
        \fpga_data_receive[3]_net_1 ), .D(\fpga_shift_2[2]_net_1 ), 
        .FCI(\fpga_flag4_0_data_tmp[0] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[1] ));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_1 (.A(
        \fpga_shift_2[1]_net_1 ), .B(\fpga_data_receive[0]_net_1 ), .C(
        \fpga_data_receive[1]_net_1 ), .D(\fpga_shift_2[0]_net_1 ), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(\fpga_flag4_0_data_tmp[0] ));
    SLE \temp_count[12]  (.D(\temp_count_s[12] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[12]));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_13 (.A(freq_6), .B(
        temp_count[13]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_12_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_13_net_1));
    CFG4 #( .INIT(16'h8000) )  temp1_14_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_178), .Y(temp1_14));
    SLE \fpga_shift[7]  (.D(\fpga_count[7]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[7]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6O6JH1[24]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[24]), .D(GND_net_1), .FCI(\temp_count_cry[23] ), .S(
        \temp_count_s[24] ), .Y(), .FCO(\temp_count_cry[24] ));
    CFG4 #( .INIT(16'h0010) )  temp2_39_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_76), .Y(temp2_39));
    CFG4 #( .INIT(16'h1000) )  temp1_26_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_178), .Y(temp1_26));
    SLE \temp_count[0]  (.D(\temp_count_s[0] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[0]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[4]  (.A(VCC_net_1), .B(
        \fpga_count[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[3]_net_1 ), .S(\fpga_count_s[4] ), .Y(), .FCO(
        \fpga_count_cry[4]_net_1 ));
    CFG3 #( .INIT(8'h94) )  \temp_state_RNIU6MV[0]  (.A(
        \temp_state[1]_net_1 ), .B(\temp_state[2]_net_1 ), .C(
        \temp_state[0]_net_1 ), .Y(N_17_i_0));
    SLE \temp1[15]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_26), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[15]));
    SLE \dac_count[8]  (.D(\dac_count_s[8]_net_1 ), .CLK(BW_clk_c), 
        .EN(clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[12]  (.A(VCC_net_1), .B(
        \cnt_freq[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[11]_net_1 ), .S(\cnt_freq_s[12] ), .Y(), .FCO(
        \cnt_freq_cry[12]_net_1 ));
    CFG4 #( .INIT(16'h3733) )  \un1_data_from_adc[2]_1lto11  (.A(
        \data_from_adc[2][9]_net_1 ), .B(\data_from_adc[2][11]_net_1 ), 
        .C(\data_from_adc[2][10]_net_1 ), .D(
        \un1_data_from_adc[2]_1lt10 ), .Y(\un1_data_from_adc[2]_1 ));
    CFG4 #( .INIT(16'h4000) )  temp2_37_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_181), .Y(temp2_37));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_4_166_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[4]_net_1 ), .Y(N_698_i));
    SLE \freq[9]  (.D(\un1_data_from_adc[2]_1_i_0 ), .CLK(temp_sck_c), 
        .EN(N_575_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(freq_2));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[8]  (.A(N_99), .B(
        \data_from_adc[2]_66_0_0_a2_0_0 ), .C(N_109), .Y(
        \data_from_adc[2]_67 ));
    SLE \temp_count[17]  (.D(\temp_count_s[17] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[17]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[6]  (.A(N_99), .B(
        \data_from_adc[2]_65_0_0_a2_1 ), .C(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .Y(\data_from_adc[2]_65 ));
    SLE \cnt_freq[7]  (.D(\cnt_freq_s[7] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[7]_net_1 ));
    SLE \fpga_shift[4]  (.D(\fpga_count[4]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[4]));
    SLE \fpga_count[3]  (.D(\fpga_count_s[3] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[3]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6US111[15]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[15]), .D(GND_net_1), .FCI(\temp_count_cry[14] ), .S(
        \temp_count_s[15] ), .Y(), .FCO(\temp_count_cry[15] ));
    SLE \temp3[12]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_55), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[12]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[17]  (.A(VCC_net_1), .B(
        \cnt_freq[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[16]_net_1 ), .S(\cnt_freq_s[17] ), .Y(), .FCO(
        \cnt_freq_cry[17]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_16 (.A(freq_1), .B(
        \cnt_freq[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_15_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_16_net_1));
    CFG4 #( .INIT(16'h82BD) )  \temp_state_7_2_0_.N_22_i  (.A(
        \temp_state[0]_net_1 ), .B(\temp_state[2]_net_1 ), .C(N_22_i_1)
        , .D(\temp_state[1]_net_1 ), .Y(N_22_i_0));
    CFG4 #( .INIT(16'h2000) )  temp2_32_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_181), .Y(temp2_32));
    SLE \data_from_adc[2][3]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_62 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][3]_net_1 ));
    SLE \cnt[3]  (.D(\cnt_s[3] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[3]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_25 (.A(VCC_net_1), .B(
        \cnt_freq[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_24_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_25_net_1));
    SLE \fpga_data_receive[1]  (.D(BW_c[1]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[1]  (.A(
        \data_from_adc[2]_68_0_0_a2_0 ), .B(N_99), .C(
        \data_from_adc[2]_66_0_0_a2_0_out ), .D(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .Y(\data_from_adc[2]_60 ));
    SLE \data_from_adc[2][10]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_69 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][10]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI7THTD1[22]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[22]), .D(GND_net_1), .FCI(\temp_count_cry[21] ), .S(
        \temp_count_s[22] ), .Y(), .FCO(\temp_count_cry[22] ));
    SLE \temp_count[1]  (.D(\temp_count_s[1] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[1]));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_8 (.A(freq_1), .B(
        temp_count[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_7_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_8_net_1));
    SLE \temp_count[20]  (.D(\temp_count_s[20] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[20]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_29 (.A(VCC_net_1), .B(
        \cnt_freq[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_28_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_29_net_1));
    SLE \temp_count[19]  (.D(\temp_count_s[19] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[19]));
    CFG4 #( .INIT(16'h0C09) )  \cnt_frame_r[2]  (.A(N_58), .B(
        \cnt_frame[2]_net_1 ), .C(cnt_frame_0_sqmuxa), .D(N_44), .Y(
        cnt_frame));
    SLE \temp_count[21]  (.D(\temp_count_s[21] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[21]));
    SLE \temp2[12]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_39), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[12]));
    CFG3 #( .INIT(8'h41) )  \cnt_frame_r[0]  (.A(cnt_frame_0_sqmuxa), 
        .B(\cnt_frame[0]_net_1 ), .C(N_44), .Y(cnt_frame_1));
    SLE \cnt[4]  (.D(\cnt_s[4] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[4]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  temp1_24_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_179), .Y(temp1_24));
    SLE \freq[22]  (.D(\un1_data_from_adc[2]_i_0 ), .CLK(temp_sck_c), 
        .EN(N_575_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(freq_15));
    SLE \cnt_freq[11]  (.D(\cnt_freq_s[11] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[11]_net_1 ));
    SLE \fpga_count[10]  (.D(\fpga_count_s[10] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[10]_net_1 ));
    SLE \temp3[3]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_46), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[3]));
    CFG4 #( .INIT(16'h6996) )  GPIO3_9 (.A(adc_d0_c[9]), .B(
        adc_d0_c[8]), .C(adc_d0_c[7]), .D(adc_d0_c[6]), .Y(
        GPIO3_9_net_1));
    SLE \dac1_db[12]  (.D(N_677_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[12]));
    SLE \cnt_freq[13]  (.D(\cnt_freq_s[13] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[13]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \cnt_RNIN2FE_0[3]  (.A(\cnt[4]_net_1 ), .B(
        \cnt[3]_net_1 ), .Y(\data_from_adc[2]_68_0_0_a2_0_out ));
    CFG3 #( .INIT(8'h80) )  \cnt_RNIBCML[1]  (.A(\cnt[2]_net_1 ), .B(
        GPIO7_c), .C(\cnt[1]_net_1 ), .Y(
        \data_from_adc[2]_68_0_0_a2_0 ));
    ARI1 #( .INIT(20'h4AAA2) )  \temp_count_RNIEEE23[0]  (.A(
        temp_count6), .B(temp_count[0]), .C(\temp_state[1]_net_1 ), .D(
        \temp_state[2]_net_1 ), .FCI(temp_count_net_1), .S(
        \temp_count_s[0] ), .Y(), .FCO(\temp_count_cry[0] ));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_5_155_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[5]_net_1 ), .Y(N_691_i));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIV5TMF[6]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[6]), .D(
        GND_net_1), .FCI(\temp_count_cry[5] ), .S(\temp_count_s[6] ), 
        .Y(), .FCO(\temp_count_cry[6] ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI771EJ1[25]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[25]), .D(GND_net_1), .FCI(\temp_count_cry[24] ), .S(
        \temp_count_s[25] ), .Y(), .FCO(\temp_count_cry[25] ));
    SLE \temp1[0]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_11), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[0]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_20 (.A(freq_13), .B(
        \cnt_freq[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_19_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_20_net_1));
    CFG4 #( .INIT(16'h4000) )  temp3_50_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_178), .Y(temp3_50));
    CFG4 #( .INIT(16'h0080) )  temp3_43_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_76), .Y(temp3_43));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[2]  (.A(VCC_net_1), .B(
        \dac_count[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[1]_net_1 ), .S(\dac_count_s[2] ), .Y(), .FCO(
        \dac_count_cry[2]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  temp1_15_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_76), .Y(temp1_15));
    CFG4 #( .INIT(16'h6996) )  GPIO5_13 (.A(osc_vcc_c), .B(adc_of_c), 
        .C(adc_oen_c), .D(adc_clk_c), .Y(GPIO5_13_net_1));
    CFG4 #( .INIT(16'h0040) )  temp2_31_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_76), .Y(temp2_31));
    SLE \fpga_count[9]  (.D(\fpga_count_s[9] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[9]_net_1 ));
    SLE \cnt_freq[28]  (.D(\cnt_freq_s[28] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[28]_net_1 ));
    CFG4 #( .INIT(16'h0020) )  temp2_csn_1_sqmuxa_0_a3 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(
        temp2_csn_1_sqmuxa));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[7]  (.A(VCC_net_1), .B(
        \fpga_count[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[6]_net_1 ), .S(\fpga_count_s[7] ), .Y(), .FCO(
        \fpga_count_cry[7]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI7CMS21[16]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[16]), .D(GND_net_1), .FCI(\temp_count_cry[15] ), .S(
        \temp_count_s[16] ), .Y(), .FCO(\temp_count_cry[16] ));
    CFG4 #( .INIT(16'h8000) )  temp2_29_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_181), .Y(temp2_29));
    SLE \data_from_adc[2][5]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_64 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][5]_net_1 ));
    SLE \dac1_db[6]  (.D(N_719_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[6]));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_12 (.A(freq_2), .B(
        \cnt_freq[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_11_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_12_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNICGNMP[11]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[11]), .D(GND_net_1), .FCI(\temp_count_cry[10] ), .S(
        \temp_count_s[11] ), .Y(), .FCO(\temp_count_cry[11] ));
    CFG4 #( .INIT(16'h51FF) )  freq15_i_0 (.A(
        \data_from_adc[2][11]_net_1 ), .B(\data_from_adc[2][10]_net_1 )
        , .C(\un1_data_from_adc[2]lt10 ), .D(\un1_data_from_adc[2]_1 ), 
        .Y(freq15_i_0_net_1));
    SLE \cnt_freq[24]  (.D(\cnt_freq_s[24] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[24]_net_1 ));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_21 (.A(
        \fpga_shift_2[9]_net_1 ), .B(\fpga_data_receive[8]_net_1 ), .C(
        \fpga_data_receive[9]_net_1 ), .D(\fpga_shift_2[8]_net_1 ), 
        .FCI(\fpga_flag4_0_data_tmp[3] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[4] ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_7 (.A(freq_0), .B(
        temp_count[7]), .C(GND_net_1), .D(GND_net_1), .FCI(GND_net_1), 
        .S(), .Y(), .FCO(temp_count6_cry_7_net_1));
    SLE \fpga_count[6]  (.D(\fpga_count_s[6] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[6]_net_1 ));
    SLE \cnt_freq[22]  (.D(\cnt_freq_s[22] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[22]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_9 (.A(freq_2), .B(
        temp_count[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_8_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_9_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[5]  (.A(VCC_net_1), .B(
        \fpga_count[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[4]_net_1 ), .S(\fpga_count_s[5] ), .Y(), .FCO(
        \fpga_count_cry[5]_net_1 ));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_0_210_x2 (.A(\sdv_count[1]_net_1 )
        , .B(GPIO20_c), .Y(N_726_i));
    CFG4 #( .INIT(16'h0080) )  temp2_27_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_76), .Y(temp2_27));
    SLE \fpga_shift_2[13]  (.D(BW_out_c[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[13]_net_1 ));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_33 (.A(
        \fpga_shift_2[5]_net_1 ), .B(\fpga_data_receive[4]_net_1 ), .C(
        \fpga_data_receive[5]_net_1 ), .D(\fpga_shift_2[4]_net_1 ), 
        .FCI(\fpga_flag4_0_data_tmp[1] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[2] ));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[2]  (.A(VCC_net_1), .B(
        N_36_i_0), .C(\cnt[2]_net_1 ), .D(GND_net_1), .FCI(
        \cnt_cry[1]_net_1 ), .S(\cnt_s[2] ), .Y(), .FCO(
        \cnt_cry[2]_net_1 ));
    SLE \temp_state[0]  (.D(N_22_i_0), .CLK(temp_sck_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_state[0]_net_1 ));
    CFG3 #( .INIT(8'h0E) )  \SENSE_DOUT_2_1_u_i_a2_0_1[1]  (.A(
        \cnt_frame[1]_net_1 ), .B(\cnt_frame[0]_net_1 ), .C(
        \cnt[2]_net_1 ), .Y(\SENSE_DOUT_2_1_u_i_a2_0_0[1]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  
        \un1_data_from_adc[2]_2lto11_i_a2_5_RNI7H6H  (.A(
        \un1_data_from_adc[2]_2lto11_i_a2_7_net_1 ), .B(
        \un1_data_from_adc[2]_2lto11_i_a2_6_net_1 ), .C(
        \un1_data_from_adc[2]_2lto11_i_a2_5_net_1 ), .Y(N_575_i_0));
    CFG4 #( .INIT(16'h8000) )  temp3_46_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_178), .Y(temp3_46));
    SLE \temp_state[2]  (.D(\temp_state_7[2] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\temp_state[2]_net_1 ));
    SLE \cnt[5]  (.D(\cnt_s[5]_net_1 ), .CLK(temp_sck_c_i_0), .EN(cnte)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[5]_net_1 ));
    SLE \fpga_shift[10]  (.D(\fpga_count[10]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[10]));
    SLE \fpga_data_receive[12]  (.D(BW_c[12]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[12]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_28 (.A(VCC_net_1), .B(
        \cnt_freq[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_27_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_28_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[24]  (.A(VCC_net_1), .B(
        \cnt_freq[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[23]_net_1 ), .S(\cnt_freq_s[24] ), .Y(), .FCO(
        \cnt_freq_cry[24]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  temp3_53_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_180), .Y(temp3_53));
    SLE \temp_count[15]  (.D(\temp_count_s[15] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[15]));
    SLE \fpga_shift[13]  (.D(\fpga_count[13]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[13]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[10]  (.A(VCC_net_1), .B(
        \cnt_freq[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[9]_net_1 ), .S(\cnt_freq_s[10] ), .Y(), .FCO(
        \cnt_freq_cry[10]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  un1_cnt_frame_0_sqmuxa_i_o4 (.A(
        \cnt[5]_net_1 ), .B(\cnt[4]_net_1 ), .C(N_54), .Y(N_52));
    CFG3 #( .INIT(8'h01) )  \SENSE_DOUT_2_1_u_i_a2_4[1]  (.A(
        \cnt_frame[3]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(
        \cnt_frame[0]_net_1 ), .Y(N_99));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[19]  (.A(VCC_net_1), .B(
        \cnt_freq[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[18]_net_1 ), .S(\cnt_freq_s[19] ), .Y(), .FCO(
        \cnt_freq_cry[19]_net_1 ));
    SLE \cnt[1]  (.D(\cnt_s[1] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[1]_net_1 ));
    SLE \fpga_shift[3]  (.D(\fpga_count[3]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[3]));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_22 (.A(freq_15), .B(
        temp_count[22]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_21_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_22_net_1));
    SLE \temp1[9]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_20), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[9]));
    CFG4 #( .INIT(16'h000D) )  \SENSE_DOUT_1_RNO[1]  (.A(N_99), .B(
        \cnt_frame[1]_net_1 ), .C(\SENSE_DOUT_2_1_u_i_1[1]_net_1 ), .D(
        N_80), .Y(N_19_i_0));
    SLE \temp3[14]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_57), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[14]));
    CFG4 #( .INIT(16'h6996) )  GPIO3_7 (.A(adc_d0_c[3]), .B(
        adc_d0_c[2]), .C(adc_d0_c[1]), .D(adc_d0_c[0]), .Y(
        GPIO3_7_net_1));
    CFG3 #( .INIT(8'h41) )  \temp_count_data_RNO[2]  (.A(
        temp_count_data[4]), .B(temp_count_data[2]), .C(N_76), .Y(
        N_10_i_0));
    SLE \fpga_count[1]  (.D(\fpga_count_s[1] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[1]_net_1 ));
    CFG2 #( .INIT(4'hE) )  temp3_csn_RNO (.A(temp_state26), .B(
        un1_temp_state_7_or), .Y(temp3_csn_RNO_net_1));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[5]  (.A(N_99), .B(
        \data_from_adc[2]_64_0_0_a2_1 ), .C(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .Y(\data_from_adc[2]_64 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[7]  (.A(VCC_net_1), .B(
        \cnt_freq[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[6]_net_1 ), .S(\cnt_freq_s[7] ), .Y(), .FCO(
        \cnt_freq_cry[7]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_17 (.A(freq_10), .B(
        temp_count[17]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_16_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_17_net_1));
    SLE \fpga_shift_2[0]  (.D(BW_out_c[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[0]_net_1 ));
    SLE \fpga_data_receive[0]  (.D(BW_c[0]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[10]  (.A(VCC_net_1), 
        .B(\fpga_count[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[9]_net_1 ), .S(\fpga_count_s[10] ), .Y(), .FCO(
        \fpga_count_cry[10]_net_1 ));
    SLE \temp1[4]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_15), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[4]));
    SLE \fpga_shift_2[3]  (.D(BW_out_c[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[3]_net_1 ));
    SLE \fpga_data_receive[6]  (.D(BW_c[6]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[6]_net_1 ));
    SLE \fpga_count[13]  (.D(\fpga_count_s[13] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[13]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_17 (.A(freq_10), .B(
        \cnt_freq[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_16_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_17_net_1));
    CFG4 #( .INIT(16'h1000) )  temp3_56_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_180), .Y(temp3_56));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[13]  (.A(VCC_net_1), 
        .B(\fpga_count[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[12]_net_1 ), .S(\fpga_count_s[13] ), .Y(), 
        .FCO(\fpga_count_cry[13]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  temp1_25_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_179), .Y(temp1_25));
    SLE \fpga_count[5]  (.D(\fpga_count_s[5] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  temp1_17_0_0_a2 (.A(temp_count_data[0]), .B(
        temp_count_data[1]), .Y(N_182));
    SLE \temp_count[5]  (.D(\temp_count_s[5] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[5]));
    SLE \temp_count[14]  (.D(\temp_count_s[14] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[14]));
    SLE \fpga_shift_2[4]  (.D(BW_out_c[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[4]_net_1 ));
    SLE \temp_count[9]  (.D(\temp_count_s[9] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[9]));
    SLE \temp3[5]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_48), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[5]));
    SLE \temp2[14]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_41), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[14]));
    SLE \fpga_shift[0]  (.D(\fpga_count[0]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[0]));
    SLE \fpga_count[7]  (.D(\fpga_count_s[7] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[7]_net_1 ));
    SLE \cnt_freq[5]  (.D(\cnt_freq_s[5] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[8]  (.A(VCC_net_1), .B(
        \cnt_freq[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[7]_net_1 ), .S(\cnt_freq_s[8] ), .Y(), .FCO(
        \cnt_freq_cry[8]_net_1 ));
    CFG3 #( .INIT(8'h01) )  SENSE_DOUT61_i_a4 (.A(\cnt[2]_net_1 ), .B(
        GPIO7_c), .C(\cnt[1]_net_1 ), .Y(N_109));
    SLE \fpga_data_receive[8]  (.D(BW_c[8]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[8]_net_1 ));
    CFG2 #( .INIT(4'h7) )  temp_count_data_n3_i_o2 (.A(
        temp_count_data[0]), .B(temp_count_data[1]), .Y(N_76));
    CFG4 #( .INIT(16'h8000) )  temp3_44_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_180), .Y(temp3_44));
    SLE \temp1[5]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_16), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[5]));
    CFG2 #( .INIT(4'hD) )  \freq_RNO[21]  (.A(\un1_data_from_adc[2]_1 )
        , .B(freq3), .Y(N_445_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[1]  (.A(VCC_net_1), .B(
        \dac_count[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        dac_count_s_460_FCO), .S(\dac_count_s[1] ), .Y(), .FCO(
        \dac_count_cry[1]_net_1 ));
    SLE \temp3[7]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_50), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[7]));
    SLE \temp3[2]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_45), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[2]));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_9 (.A(
        \fpga_shift_2[13]_net_1 ), .B(\fpga_data_receive[12]_net_1 ), 
        .C(\fpga_data_receive[13]_net_1 ), .D(\fpga_shift_2[12]_net_1 )
        , .FCI(\fpga_flag4_0_data_tmp[5] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[6] ));
    SLE \data_from_adc[2][8]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_67 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][8]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_9 (.A(freq_2), .B(
        \cnt_freq[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_8_net_1), .S(), .Y(), .FCO(cnt_freq6_cry_9_net_1)
        );
    SLE \cnt_freq[31]  (.D(\cnt_freq_s[31]_net_1 ), .CLK(temp_sck_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        cnt_freq6), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \cnt_freq[31]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIG7URN[10]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[10]), .D(GND_net_1), .FCI(\temp_count_cry[9] ), .S(
        \temp_count_s[10] ), .Y(), .FCO(\temp_count_cry[10] ));
    CFG4 #( .INIT(16'h6996) )  GPIO5_12 (.A(GPIO6_c), .B(GPIO4_c), .C(
        ANTF_n2_c), .D(ANTF_n1_c), .Y(GPIO5_12_net_1));
    CFG2 #( .INIT(4'h4) )  \cnt_RNIN2FE[3]  (.A(\cnt[4]_net_1 ), .B(
        \cnt[3]_net_1 ), .Y(\data_from_adc[2]_66_0_0_a2_0_out ));
    SLE \fpga_shift[6]  (.D(\fpga_count[6]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[6]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[3]  (.A(VCC_net_1), .B(
        \cnt_freq[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[2]_net_1 ), .S(\cnt_freq_s[3] ), .Y(), .FCO(
        \cnt_freq_cry[3]_net_1 ));
    CFG4 #( .INIT(16'h010A) )  \state_RNO[1]  (.A(\state[1]_net_1 ), 
        .B(\cnt_frame[3]_net_1 ), .C(N_86), .D(\state[0]_net_1 ), .Y(
        N_23_i_0));
    SLE \fpga_data_receive[3]  (.D(BW_c[3]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[3]_net_1 ));
    SLE \temp3[13]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_56), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[13]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_23 (.A(VCC_net_1), .B(
        \cnt_freq[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_22_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_23_net_1));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_21 (.A(freq_14), .B(
        \cnt_freq[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_20_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_21_net_1));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_14 (.A(VCC_net_1), .B(
        temp_count[14]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_13_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_14_net_1));
    SLE \fpga_shift[1]  (.D(\fpga_count[1]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[1]));
    SLE \fpga_data_receive[5]  (.D(BW_c[5]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[5]_net_1 ));
    CFG4 #( .INIT(16'h4451) )  temp1_csn_RNO_0 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(
        un1_temp_state_8_or));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[12]  (.A(VCC_net_1), 
        .B(\fpga_count[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[11]_net_1 ), .S(\fpga_count_s[12] ), .Y(), 
        .FCO(\fpga_count_cry[12]_net_1 ));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_3_177_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[3]_net_1 ), .Y(N_705_i));
    SLE temp3_csn (.D(\temp_state[1]_net_1 ), .CLK(temp_sck_c), .EN(
        temp3_csn_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_322_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(temp3_csn_c));
    SLE temp1_csn (.D(\temp_state[0]_net_1 ), .CLK(temp_sck_c), .EN(
        temp1_csn_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_322_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(temp1_csn_c));
    SLE \cnt_freq[19]  (.D(\cnt_freq_s[19] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[19]_net_1 ));
    CFG4 #( .INIT(16'hC8CC) )  \un1_data_from_adc[2]_1lto11_i  (.A(
        \data_from_adc[2][9]_net_1 ), .B(\data_from_adc[2][11]_net_1 ), 
        .C(\data_from_adc[2][10]_net_1 ), .D(
        \un1_data_from_adc[2]_1lt10 ), .Y(\un1_data_from_adc[2]_1_i_0 )
        );
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_29 (.A(VCC_net_1), .B(
        temp_count[29]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_28_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_29_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[23]  (.A(VCC_net_1), .B(
        \cnt_freq[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[22]_net_1 ), .S(\cnt_freq_s[23] ), .Y(), .FCO(
        \cnt_freq_cry[23]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_1_199_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[1]_net_1 ), .Y(N_719_i));
    SLE \temp3[15]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_58), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[15]));
    CFG4 #( .INIT(16'h2000) )  temp2_38_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_178), .Y(temp2_38));
    CFG4 #( .INIT(16'hFEFF) )  freq3lto11_i (.A(
        \data_from_adc[2][9]_net_1 ), .B(\data_from_adc[2][11]_net_1 ), 
        .C(\data_from_adc[2][10]_net_1 ), .D(freq3lt11), .Y(freq3_i_0));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_27 (.A(
        \fpga_shift_2[7]_net_1 ), .B(\fpga_data_receive[6]_net_1 ), .C(
        \fpga_data_receive[7]_net_1 ), .D(\fpga_shift_2[6]_net_1 ), 
        .FCI(\fpga_flag4_0_data_tmp[2] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[3] ));
    SLE \dac1_db[5]  (.D(N_726_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[5]));
    CFG1 #( .INIT(2'h1) )  \temp_state_RNI91IA[0]  (.A(
        \temp_state[0]_net_1 ), .Y(\temp_state_i_0[0] ));
    CFG4 #( .INIT(16'h2000) )  temp3_54_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_178), .Y(temp3_54));
    CFG2 #( .INIT(4'h7) )  \state_RNI9IAG[1]  (.A(\state[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(N_70_i_0));
    CFG4 #( .INIT(16'h6996) )  GPIO3_8 (.A(adc_d0_c[13]), .B(
        adc_d0_c[12]), .C(adc_d0_c[11]), .D(adc_d0_c[10]), .Y(
        GPIO3_8_net_1));
    SLE \temp2[13]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_40), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[13]));
    SLE \cnt_freq[4]  (.D(\cnt_freq_s[4] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[4]_net_1 ));
    SLE \fpga_shift_2[6]  (.D(BW_out_c[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[6]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_24 (.A(VCC_net_1), .B(
        \cnt_freq[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_23_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_24_net_1));
    CFG3 #( .INIT(8'h7F) )  \un1_data_from_adc[2]lto4  (.A(
        \data_from_adc[2][2]_net_1 ), .B(\data_from_adc[2][4]_net_1 ), 
        .C(\data_from_adc[2][3]_net_1 ), .Y(\un1_data_from_adc[2]lt5 ));
    CFG4 #( .INIT(16'h0004) )  temp1_11_0_0_a2 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(N_179));
    CFG2 #( .INIT(4'h1) )  freq3lto3 (.A(\data_from_adc[2][2]_net_1 ), 
        .B(\data_from_adc[2][3]_net_1 ), .Y(freq3lt8));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[4]  (.A(VCC_net_1), .B(
        \cnt_freq[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[3]_net_1 ), .S(\cnt_freq_s[4] ), .Y(), .FCO(
        \cnt_freq_cry[4]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \SENSE_DOUT_2_1_u_i_a2_0[1]  (.A(N_58), 
        .B(\SENSE_DOUT_2_1_u_i_a2_0_0[1]_net_1 ), .C(\cnt[1]_net_1 ), 
        .D(GPIO7_c), .Y(N_43));
    CFG3 #( .INIT(8'h46) )  \SENSE_DOUT_2_1_u_i_1_RNO[1]  (.A(
        \cnt_frame[2]_net_1 ), .B(\cnt_frame[1]_net_1 ), .C(
        \cnt_frame[0]_net_1 ), .Y(N_3563_tz));
    SLE \cnt_freq[3]  (.D(\cnt_freq_s[3] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[3]_net_1 ));
    SLE \temp_count[28]  (.D(\temp_count_s[28] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[28]));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_31 (.A(VCC_net_1), .B(
        temp_count[31]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_30_net_1), .S(), .Y(), .FCO(temp_count6));
    CFG4 #( .INIT(16'h6620) )  temp2_csn_RNO_0 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(
        un1_temp_state29_3_or));
    SLE \temp2[15]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_42), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[15]));
    CFG4 #( .INIT(16'hF1F0) )  \un1_data_from_adc[2]_1lto8  (.A(
        \data_from_adc[2][4]_net_1 ), .B(\data_from_adc[2][5]_net_1 ), 
        .C(\un1_data_from_adc[2]lto8_0_net_1 ), .D(freq3lt8), .Y(
        \un1_data_from_adc[2]_1lt10 ));
    SLE \temp2[8]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_35), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[8]));
    CFG2 #( .INIT(4'h4) )  SENSE_CS_1_RNIM4KA (.A(SENSE_CS_1_c), .B(
        temp_sck_c), .Y(oclk_1_c));
    CFG3 #( .INIT(8'hF2) )  \freq_RNO[22]  (.A(
        \data_from_adc[2][10]_net_1 ), .B(\un1_data_from_adc[2]lt10 ), 
        .C(\data_from_adc[2][11]_net_1 ), .Y(
        \un1_data_from_adc[2]_i_0 ));
    CFG4 #( .INIT(16'hF1FA) )  \cnt_frame_RNI0N272[3]  (.A(
        \state[1]_net_1 ), .B(\cnt_frame[3]_net_1 ), .C(N_36_i_0), .D(
        \state[0]_net_1 ), .Y(cnte));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_16 (.A(freq_1), .B(
        temp_count[16]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_15_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_16_net_1));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_25 (.A(VCC_net_1), .B(
        temp_count[25]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_24_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_25_net_1));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI0Q2GB[4]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[4]), .D(
        GND_net_1), .FCI(\temp_count_cry[3] ), .S(\temp_count_s[4] ), 
        .Y(), .FCO(\temp_count_cry[4] ));
    CFG4 #( .INIT(16'h4414) )  \temp_count_data_RNO[3]  (.A(
        temp_count_data[4]), .B(temp_count_data[3]), .C(
        temp_count_data[2]), .D(N_76), .Y(N_8_i_0));
    CFG4 #( .INIT(16'h0020) )  temp1_19_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_76), .Y(temp1_19));
    SLE \fpga_data_receive[13]  (.D(BW_c[13]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[13]_net_1 ));
    SLE \fpga_shift[12]  (.D(\fpga_count[12]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[12]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_30 (.A(VCC_net_1), .B(
        \cnt_freq[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_29_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_30_net_1));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[3]  (.A(VCC_net_1), .B(
        N_36_i_0), .C(\cnt[3]_net_1 ), .D(GND_net_1), .FCI(
        \cnt_cry[2]_net_1 ), .S(\cnt_s[3] ), .Y(), .FCO(
        \cnt_cry[3]_net_1 ));
    SLE \temp_count[8]  (.D(\temp_count_s[8] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[8]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI5I897[2]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[2]), .D(
        GND_net_1), .FCI(\temp_count_cry[1] ), .S(\temp_count_s[2] ), 
        .Y(), .FCO(\temp_count_cry[2] ));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[0]  (.A(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .B(
        \data_from_adc[2]_59_0_0_a2_0 ), .C(N_99), .D(N_109), .Y(
        \data_from_adc[2]_59 ));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_2_188_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[2]_net_1 ), .Y(N_712_i));
    SLE \cnt_frame[2]  (.D(cnt_frame), .CLK(temp_sck_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_frame[2]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \cnt_cry[0]  (.A(VCC_net_1), .B(
        GPIO7_c), .C(N_36_i_0), .D(GND_net_1), .FCI(cnt_cry_cy), .S(
        \cnt_s[0] ), .Y(), .FCO(\cnt_cry[0]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIC6T7A1[20]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[20]), .D(GND_net_1), .FCI(\temp_count_cry[19] ), .S(
        \temp_count_s[20] ), .Y(), .FCO(\temp_count_cry[20] ));
    CFG3 #( .INIT(8'h02) )  \data_from_adc[2]_RNO_0[4]  (.A(
        \cnt[2]_net_1 ), .B(GPIO7_c), .C(\cnt[1]_net_1 ), .Y(
        \data_from_adc[2]_63_0_0_a2_0 ));
    ARI1 #( .INIT(20'h49900) )  fpga_flag4_0_I_45 (.A(VCC_net_1), .B(
        \fpga_data_receive[14]_net_1 ), .C(\fpga_shift_2[14]_net_1 ), 
        .D(GND_net_1), .FCI(\fpga_flag4_0_data_tmp[6] ), .S(), .Y(), 
        .FCO(fpga_flags));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_s[31]  (.A(VCC_net_1), .B(
        \cnt_freq[31]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[30]_net_1 ), .S(\cnt_freq_s[31]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_20 (.A(freq_13), .B(
        temp_count[20]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_19_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_20_net_1));
    CFG4 #( .INIT(16'h2000) )  temp1_17_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_179), .Y(temp1_17));
    SLE \fpga_shift_2[8]  (.D(BW_out_c[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[15]  (.A(VCC_net_1), .B(
        \cnt_freq[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[14]_net_1 ), .S(\cnt_freq_s[15] ), .Y(), .FCO(
        \cnt_freq_cry[15]_net_1 ));
    CFG3 #( .INIT(8'hFD) )  \cnt_frame_0_i_o4[0]  (.A(\state[0]_net_1 )
        , .B(\cnt_frame[3]_net_1 ), .C(\state[1]_net_1 ), .Y(N_44));
    CFG4 #( .INIT(16'h8000) )  temp3_45_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_180), .Y(temp3_45));
    CFG4 #( .INIT(16'h6996) )  GPIO5_11 (.A(GPS1_LD_c), .B(GPS1_I1_c), 
        .C(GPS1_I0_c), .D(GPIO9_c), .Y(GPIO5_11_net_1));
    SLE GPIO16 (.D(N_12_i_0), .CLK(temp_sck_c), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(GPIO16_c));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI2MNTJ[8]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[8]), .D(
        GND_net_1), .FCI(\temp_count_cry[7] ), .S(\temp_count_s[8] ), 
        .Y(), .FCO(\temp_count_cry[8] ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_23 (.A(VCC_net_1), .B(
        temp_count[23]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_22_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_23_net_1));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[11]  (.A(
        \data_from_adc[2]_70_0_0_a2_0 ), .B(N_99), .C(
        \data_from_adc[2]_68_0_0_a2_0_out ), .D(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .Y(\data_from_adc[2]_70 ));
    CFG4 #( .INIT(16'h0002) )  temp2_27_0_0_a2 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(N_181));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_26 (.A(VCC_net_1), .B(
        \cnt_freq[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_25_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_26_net_1));
    SLE clk_dac1 (.D(clk_dac1_2_net_1), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dac1_clk_c));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[1]  (.A(VCC_net_1), .B(
        \fpga_count[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        fpga_count_s_459_FCO), .S(\fpga_count_s[1] ), .Y(), .FCO(
        \fpga_count_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_s[14]  (.A(VCC_net_1), .B(
        \fpga_count[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[13]_net_1 ), .S(\fpga_count_s[14]_net_1 ), .Y()
        , .FCO());
    ARI1 #( .INIT(20'h4EF00) )  temp_count6_cry_31_RNIPJ5K1 (.A(
        VCC_net_1), .B(temp_count6), .C(\temp_state[2]_net_1 ), .D(
        \temp_state[1]_net_1 ), .FCI(temp_count_lcry_cy), .S(), .Y(
        temp_count6_cry_31_RNIPJ5K1_Y), .FCO(temp_count_net_1));
    SLE \temp_count[16]  (.D(\temp_count_s[16] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[16]));
    CFG3 #( .INIT(8'h20) )  \cnt_RNIBCML_0[1]  (.A(\cnt[2]_net_1 ), .B(
        GPIO7_c), .C(\cnt[1]_net_1 ), .Y(\data_from_adc[2]_61_1 ));
    SLE \temp2[4]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_31), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[4]));
    CFG4 #( .INIT(16'h8000) )  temp1_12_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_179), .Y(temp1_12));
    SLE \fpga_shift_2[12]  (.D(BW_out_c[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[30]  (.A(VCC_net_1), .B(
        \cnt_freq[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[29]_net_1 ), .S(\cnt_freq_s[30] ), .Y(), .FCO(
        \cnt_freq_cry[30]_net_1 ));
    SLE \temp_count_data[2]  (.D(N_10_i_0), .CLK(temp_sck_c), .EN(
        N_17_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count_data[2]));
    SLE \temp2[9]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_36), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[9]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[9]  (.A(VCC_net_1), .B(
        \cnt_freq[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[8]_net_1 ), .S(\cnt_freq_s[9] ), .Y(), .FCO(
        \cnt_freq_cry[9]_net_1 ));
    CFG4 #( .INIT(16'h3310) )  \un1_data_from_adc[2]lto9  (.A(
        \data_from_adc[2][5]_net_1 ), .B(\data_from_adc[2][9]_net_1 ), 
        .C(\un1_data_from_adc[2]lt5 ), .D(
        \un1_data_from_adc[2]lto8_0_net_1 ), .Y(
        \un1_data_from_adc[2]lt10 ));
    SLE \temp2[5]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_32), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[5]));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_8_122_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[8]_net_1 ), .Y(N_670_i));
    CFG4 #( .INIT(16'h8000) )  temp2_28_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_181), .Y(temp2_28));
    SLE \fpga_data_receive[11]  (.D(BW_c[11]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[11]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \un1_data_from_adc[2]lto8_0  (.A(
        \data_from_adc[2][8]_net_1 ), .B(\data_from_adc[2][7]_net_1 ), 
        .C(\data_from_adc[2][6]_net_1 ), .Y(
        \un1_data_from_adc[2]lto8_0_net_1 ));
    SLE \dac_count[7]  (.D(\dac_count_s[7] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[7]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[3]  (.A(VCC_net_1), .B(
        \fpga_count[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[2]_net_1 ), .S(\fpga_count_s[3] ), .Y(), .FCO(
        \fpga_count_cry[3]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  temp3_55_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_76), .Y(temp3_55));
    CFG4 #( .INIT(16'h8000) )  temp2_30_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_178), .Y(temp2_30));
    SLE \sdv_count[1]  (.D(\sdv_count_1[1] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\sdv_count[1]_net_1 ));
    SLE \fpga_shift_2[1]  (.D(BW_out_c[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[4]  (.A(VCC_net_1), .B(
        \dac_count[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[3]_net_1 ), .S(\dac_count_s[4] ), .Y(), .FCO(
        \dac_count_cry[4]_net_1 ));
    SLE clk_dac2 (.D(\sdv_count[0]_net_1 ), .CLK(BW_clk_c), .EN(
        \sdv_count[1]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(clk_dac2_net_1)
        );
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNO[31]  (.A(VCC_net_1), 
        .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[31]), .D(
        GND_net_1), .FCI(\temp_count_cry[30] ), .S(\temp_count_s[31] ), 
        .Y(), .FCO());
    CFG2 #( .INIT(4'hE) )  \cnt_frame_RNO[3]  (.A(
        \cnt_frame_0_0_a2_0_2[3]_net_1 ), .B(cnt_frame_0_sqmuxa), .Y(
        \cnt_frame_RNO[3]_net_1 ));
    SLE \cnt_freq[9]  (.D(\cnt_freq_s[9] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[9]_net_1 ));
    SLE \temp_count[2]  (.D(\temp_count_s[2] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[2]));
    SLE \temp_count[22]  (.D(\temp_count_s[22] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[22]));
    SLE \data_from_adc[2][9]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_68 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][9]_net_1 ));
    SLE \SENSE_DOUT_1[1]  (.D(N_19_i_0), .CLK(temp_sck_c_i_0), .EN(
        N_39_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(SENSE_DOUT_c[1]));
    CFG4 #( .INIT(16'h110A) )  un1_cnt_frame_0_sqmuxa_i_o4_RNIIAS91 (
        .A(\state[1]_net_1 ), .B(\cnt_frame[3]_net_1 ), .C(N_52), .D(
        \state[0]_net_1 ), .Y(N_36_i_0));
    CFG3 #( .INIT(8'h20) )  temp_state26_0_a3 (.A(
        \temp_state[1]_net_1 ), .B(\temp_state[2]_net_1 ), .C(
        \temp_state[0]_net_1 ), .Y(temp_state26));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIFVFJD[5]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[5]), .D(
        GND_net_1), .FCI(\temp_count_cry[4] ), .S(\temp_count_s[5] ), 
        .Y(), .FCO(\temp_count_cry[5] ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[28]  (.A(VCC_net_1), .B(
        \cnt_freq[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[27]_net_1 ), .S(\cnt_freq_s[28] ), .Y(), .FCO(
        \cnt_freq_cry[28]_net_1 ));
    SLE \fpga_shift[9]  (.D(\fpga_count[9]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[9]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[26]  (.A(VCC_net_1), .B(
        \cnt_freq[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[25]_net_1 ), .S(\cnt_freq_s[26] ), .Y(), .FCO(
        \cnt_freq_cry[26]_net_1 ));
    SLE \temp_count_data[0]  (.D(N_113), .CLK(temp_sck_c), .EN(
        N_17_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count_data[0]));
    SLE \temp_count[4]  (.D(\temp_count_s[4] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[4]));
    SLE \fpga_shift_2[5]  (.D(BW_out_c[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[5]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_22 (.A(freq_15), .B(
        \cnt_freq[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_21_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_22_net_1));
    SLE \temp_count[13]  (.D(\temp_count_s[13] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[13]));
    SLE \temp1[6]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_17), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[6]));
    CFG4 #( .INIT(16'h0080) )  temp1_11_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_76), .Y(temp1_11));
    SLE \cnt_freq[15]  (.D(\cnt_freq_s[15] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[15]_net_1 ));
    SLE \fpga_shift_2[9]  (.D(BW_out_c[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[9]_net_1 ));
    SLE \fpga_shift[2]  (.D(\fpga_count[2]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[2]));
    SLE \cnt_freq[21]  (.D(\cnt_freq_s[21] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[21]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9RFN41[17]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[17]), .D(GND_net_1), .FCI(\temp_count_cry[16] ), .S(
        \temp_count_s[17] ), .Y(), .FCO(\temp_count_cry[17] ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6ACOF1[23]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[23]), .D(GND_net_1), .FCI(\temp_count_cry[22] ), .S(
        \temp_count_s[23] ), .Y(), .FCO(\temp_count_cry[23] ));
    SLE \temp_count[27]  (.D(\temp_count_s[27] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[27]));
    CFG4 #( .INIT(16'h1000) )  temp2_42_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_178), .Y(temp2_42));
    SLE \fpga_count[8]  (.D(\fpga_count_s[8] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[8]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \sdv_count_RNO[1]  (.A(\sdv_count[1]_net_1 )
        , .B(\sdv_count[0]_net_1 ), .Y(\sdv_count_1[1] ));
    SLE \cnt_freq[23]  (.D(\cnt_freq_s[23] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[23]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIGS2D81[19]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[19]), .D(GND_net_1), .FCI(\temp_count_cry[18] ), .S(
        \temp_count_s[19] ), .Y(), .FCO(\temp_count_cry[19] ));
    CFG4 #( .INIT(16'h2000) )  temp2_33_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_181), .Y(temp2_33));
    CFG1 #( .INIT(2'h1) )  temp_state26_0_a3_RNIBC45 (.A(temp_state26), 
        .Y(N_322_i));
    SLE \cnt_frame[0]  (.D(cnt_frame_1), .CLK(temp_sck_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_frame[0]_net_1 ));
    SLE \dac1_db[7]  (.D(N_712_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[7]));
    SLE \cnt_freq[10]  (.D(\cnt_freq_s[10] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[10]_net_1 ));
    SLE \temp_state[1]  (.D(N_11_i_0), .CLK(temp_sck_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_state[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[21]  (.A(VCC_net_1), .B(
        \cnt_freq[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[20]_net_1 ), .S(\cnt_freq_s[21] ), .Y(), .FCO(
        \cnt_freq_cry[21]_net_1 ));
    SLE \temp3[6]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_49), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[6]));
    CFG4 #( .INIT(16'h2000) )  temp1_22_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_178), .Y(temp1_22));
    SLE \dac_count[1]  (.D(\dac_count_s[1] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \cnt_freq_RNO[0]  (.A(\cnt_freq[0]_net_1 ), 
        .Y(\cnt_freq_s[0] ));
    SLE \dac1_db[10]  (.D(N_691_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[10]));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_31 (.A(VCC_net_1), .B(
        \cnt_freq[31]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_30_net_1), .S(), .Y(), .FCO(cnt_freq6));
    SLE \temp2[6]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_33), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[6]));
    SLE \cnt_freq[17]  (.D(\cnt_freq_s[17] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[17]_net_1 ));
    SLE \temp1[10]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_21), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[10]));
    SLE \fpga_shift[14]  (.D(\fpga_count[14]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[14]));
    CFG1 #( .INIT(2'h1) )  clk_dac1_2_RNO (.A(\sdv_count[1]_net_1 ), 
        .Y(\sdv_count_i_0[1] ));
    CFG4 #( .INIT(16'hCCCE) )  \SENSE_DOUT_2_1_u_i_1[1]  (.A(N_3563_tz)
        , .B(N_43), .C(\cnt[2]_net_1 ), .D(GPIO7_c), .Y(
        \SENSE_DOUT_2_1_u_i_1[1]_net_1 ));
    SLE \freq[18]  (.D(\un1_data_from_adc[2]_1 ), .CLK(temp_sck_c), 
        .EN(N_575_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(freq_11));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[11]  (.A(VCC_net_1), 
        .B(\fpga_count[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[10]_net_1 ), .S(\fpga_count_s[11] ), .Y(), 
        .FCO(\fpga_count_cry[11]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  temp2_36_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_181), .Y(temp2_36));
    CFG4 #( .INIT(16'h0040) )  \data_from_adc[2]_RNO_0[6]  (.A(GPIO7_c)
        , .B(\data_from_adc[2]_66_0_0_a2_0_out ), .C(\cnt[1]_net_1 ), 
        .D(\cnt[2]_net_1 ), .Y(\data_from_adc[2]_65_0_0_a2_1 ));
    CFG3 #( .INIT(8'h40) )  \cnt_RNINDI21[5]  (.A(\cnt[5]_net_1 ), .B(
        \cnt_frame[1]_net_1 ), .C(\data_from_adc[2]_66_0_0_a2_0_out ), 
        .Y(\data_from_adc[2]_66_0_0_a2_0_0 ));
    CFG2 #( .INIT(4'h4) )  \SENSE_DOUT_2_1_u_i_a2_0_0[1]  (.A(GPIO7_c), 
        .B(\cnt_frame[0]_net_1 ), .Y(
        \SENSE_DOUT_2_1_u_i_a2_0[1]_net_1 ));
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[4]  (.A(VCC_net_1), .B(
        N_36_i_0), .C(\cnt[4]_net_1 ), .D(GND_net_1), .FCI(
        \cnt_cry[3]_net_1 ), .S(\cnt_s[4] ), .Y(), .FCO(
        \cnt_cry[4]_net_1 ));
    SLE \temp_count[29]  (.D(\temp_count_s[29] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[29]));
    SLE \temp2[3]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_30), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[3]));
    SLE \data_from_adc[2][4]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_63 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][4]_net_1 ));
    SLE \dac_count[0]  (.D(\dac_count_s[0] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(GPIO20_c));
    ARI1 #( .INIT(20'h45500) )  cnt_freq6_cry_27 (.A(VCC_net_1), .B(
        \cnt_freq[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_26_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_27_net_1));
    CFG4 #( .INIT(16'h1000) )  temp2_41_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_181), .Y(temp2_41));
    CFG2 #( .INIT(4'h8) )  clk_dac2_RNIJBB8 (.A(GPIO10_c), .B(
        clk_dac2_net_1), .Y(dac2_clk_c));
    CFG4 #( .INIT(16'h10BF) )  \temp_state_7_2_0_.N_22_i_1  (.A(
        \temp_state[2]_net_1 ), .B(GPIO11_c), .C(\temp_state[1]_net_1 )
        , .D(temp_count_data[4]), .Y(N_22_i_1));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_7 (.A(freq_0), .B(
        \cnt_freq[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(cnt_freq6_cry_7_net_1));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[7]  (.A(GPIO7_c), 
        .B(\data_from_adc[2]_66_0_0_a2_0 ), .C(N_99), .D(
        \data_from_adc[2]_66_0_0_a2_0_0 ), .Y(\data_from_adc[2]_66 ));
    ARI1 #( .INIT(20'h44400) )  \cnt_s[5]  (.A(VCC_net_1), .B(N_36_i_0)
        , .C(\cnt[5]_net_1 ), .D(GND_net_1), .FCI(\cnt_cry[4]_net_1 ), 
        .S(\cnt_s[5]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h44400) )  \cnt_cry[1]  (.A(VCC_net_1), .B(
        N_36_i_0), .C(\cnt[1]_net_1 ), .D(GND_net_1), .FCI(
        \cnt_cry[0]_net_1 ), .S(\cnt_s[1] ), .Y(), .FCO(
        \cnt_cry[1]_net_1 ));
    SLE \temp1[11]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_22), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[11]));
    SLE \freq[15]  (.D(freq9_net_1), .CLK(temp_sck_c), .EN(N_575_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(freq_0));
    SLE \cnt_freq[2]  (.D(\cnt_freq_s[2] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[2]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  GPIO5_14 (.A(GPIO5_10_net_1), .B(
        GPS_I1_c), .C(GPS_I0_c), .D(GPS2_Q1_c), .Y(GPIO5_14_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[22]  (.A(VCC_net_1), .B(
        \cnt_freq[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[21]_net_1 ), .S(\cnt_freq_s[22] ), .Y(), .FCO(
        \cnt_freq_cry[22]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_11 (.A(freq_1), .B(
        temp_count[11]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_10_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_11_net_1));
    SLE \fpga_shift[11]  (.D(\fpga_count[11]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[11]));
    SLE \dac_count[3]  (.D(\dac_count_s[3] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[3]_net_1 ));
    SLE \cnt_freq[16]  (.D(\cnt_freq_s[16] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[16]_net_1 ));
    CFG4 #( .INIT(16'hAE00) )  freq15 (.A(\data_from_adc[2][11]_net_1 )
        , .B(\data_from_adc[2][10]_net_1 ), .C(
        \un1_data_from_adc[2]lt10 ), .D(\un1_data_from_adc[2]_1 ), .Y(
        freq15_net_1));
    CFG4 #( .INIT(16'h2227) )  \temp_state_7_2_0_.m10_0_0  (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(m10_0_0));
    CFG4 #( .INIT(16'h4000) )  temp1_21_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_179), .Y(temp1_21));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[6]  (.A(VCC_net_1), .B(
        \cnt_freq[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[5]_net_1 ), .S(\cnt_freq_s[6] ), .Y(), .FCO(
        \cnt_freq_cry[6]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_18 (.A(freq_11), .B(
        temp_count[18]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_17_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_18_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[2]  (.A(VCC_net_1), .B(
        \cnt_freq[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[1]_net_1 ), .S(\cnt_freq_s[2] ), .Y(), .FCO(
        \cnt_freq_cry[2]_net_1 ));
    SLE \temp3[4]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_47), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[4]));
    CFG4 #( .INIT(16'h2AEA) )  \temp_state_7_2_0_.m13_0  (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(
        \temp_state_7[2] ));
    SLE \temp_count_data[4]  (.D(N_6_i_0), .CLK(temp_sck_c), .EN(
        N_17_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count_data[4]));
    SLE \temp1[2]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_13), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[2]));
    SLE \fpga_shift_2[14]  (.D(BW_out_c[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[14]_net_1 ));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_7_133_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[7]_net_1 ), .Y(N_677_i));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNILV41M[9]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[9]), .D(
        GND_net_1), .FCI(\temp_count_cry[8] ), .S(\temp_count_s[9] ), 
        .Y(), .FCO(\temp_count_cry[9] ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_27 (.A(VCC_net_1), .B(
        temp_count[27]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_26_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_27_net_1));
    SLE fpga_flag (.D(fpga_flags), .CLK(BW_clk_c_i_0), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(fpga_flag_i), .SD(
        VCC_net_1), .LAT(GND_net_1), .Q(fpga_flag_net_1));
    CFG2 #( .INIT(4'h6) )  dac1_db_4_6_144_x2 (.A(\sdv_count[1]_net_1 )
        , .B(\dac_count[6]_net_1 ), .Y(N_684_i));
    SLE \fpga_data_receive[10]  (.D(BW_c[10]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[10]_net_1 ));
    SLE \fpga_shift_2[2]  (.D(BW_out_c[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[14]  (.A(VCC_net_1), .B(
        \cnt_freq[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[13]_net_1 ), .S(\cnt_freq_s[14] ), .Y(), .FCO(
        \cnt_freq_cry[14]_net_1 ));
    SLE \dac_count[4]  (.D(\dac_count_s[4] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[4]_net_1 ));
    CFG3 #( .INIT(8'h01) )  cnt_frame_0_sqmuxa_0_a2 (.A(
        \state[0]_net_1 ), .B(GPIO11_c), .C(\state[1]_net_1 ), .Y(
        cnt_frame_0_sqmuxa));
    CFG4 #( .INIT(16'h2000) )  temp3_49_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_180), .Y(temp3_49));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[27]  (.A(VCC_net_1), .B(
        \cnt_freq[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[26]_net_1 ), .S(\cnt_freq_s[27] ), .Y(), .FCO(
        \cnt_freq_cry[27]_net_1 ));
    SLE \temp_count[10]  (.D(\temp_count_s[10] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[10]));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[8]  (.A(VCC_net_1), .B(
        \fpga_count[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[7]_net_1 ), .S(\fpga_count_s[8] ), .Y(), .FCO(
        \fpga_count_cry[8]_net_1 ));
    SLE \temp1[8]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_19), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[8]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIIP6KS1[30]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[30]), .D(GND_net_1), .FCI(\temp_count_cry[29] ), .S(
        \temp_count_s[30] ), .Y(), .FCO(\temp_count_cry[30] ));
    CFG2 #( .INIT(4'h2) )  \data_from_adc[2]_RNO_0[0]  (.A(
        \cnt[4]_net_1 ), .B(\cnt[3]_net_1 ), .Y(
        \data_from_adc[2]_59_0_0_a2_0 ));
    SLE \cnt_frame[3]  (.D(VCC_net_1), .CLK(temp_sck_c_i_0), .EN(
        \cnt_frame_RNO[3]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(N_333_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \cnt_frame[3]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIPFR55[1]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[1]), .D(
        GND_net_1), .FCI(\temp_count_cry[0] ), .S(\temp_count_s[1] ), 
        .Y(), .FCO(\temp_count_cry[1] ));
    SLE \temp_count[11]  (.D(\temp_count_s[11] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[11]));
    SLE \temp3[9]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_52), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[9]));
    CFG4 #( .INIT(16'h4000) )  temp2_34_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_178), .Y(temp2_34));
    CFG4 #( .INIT(16'h0040) )  temp3_47_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_76), .Y(temp3_47));
    SLE \temp1[1]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_12), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[1]));
    CFG4 #( .INIT(16'hE6EE) )  SENSE_CS_1_4_iv_i_0 (.A(\cnt[5]_net_1 ), 
        .B(\cnt[4]_net_1 ), .C(SENSE_CS_1_c), .D(N_54), .Y(N_21));
    SLE \temp_count[25]  (.D(\temp_count_s[25] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[25]));
    SLE \freq[20]  (.D(freq15_i_0_net_1), .CLK(temp_sck_c), .EN(
        N_575_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(freq_13));
    CFG4 #( .INIT(16'h0C06) )  \cnt_frame_r[1]  (.A(
        \cnt_frame[0]_net_1 ), .B(\cnt_frame[1]_net_1 ), .C(
        cnt_frame_0_sqmuxa), .D(N_44), .Y(cnt_frame_0));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[1]  (.A(VCC_net_1), .B(
        \cnt_freq[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq_s_461_FCO), .S(\cnt_freq_s[1] ), .Y(), .FCO(
        \cnt_freq_cry[1]_net_1 ));
    SLE \temp3[1]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_44), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[1]));
    SLE \temp2[1]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_28), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[1]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIC8M3N1[27]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[27]), .D(GND_net_1), .FCI(\temp_count_cry[26] ), .S(
        \temp_count_s[27] ), .Y(), .FCO(\temp_count_cry[27] ));
    SLE \cnt_freq[6]  (.D(\cnt_freq_s[6] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[6]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  temp1_18_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_179), .D(N_178), .Y(temp1_18));
    CFG1 #( .INIT(2'h1) )  \dac_count_RNO[0]  (.A(GPIO20_c), .Y(
        \dac_count_s[0] ));
    ARI1 #( .INIT(20'h42200) )  \temp_state_RNIL54L[2]  (.A(VCC_net_1), 
        .B(\temp_state[1]_net_1 ), .C(\temp_state[2]_net_1 ), .D(
        GND_net_1), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        temp_count_lcry_cy));
    CFG2 #( .INIT(4'h6) )  GPIO3_6 (.A(adc_d0_c[4]), .B(adc_d0_c[5]), 
        .Y(GPIO3_6_net_1));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[10]  (.A(
        \data_from_adc[2]_68_0_0_a2_0_out ), .B(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .C(\data_from_adc[2]_61_1 ), 
        .D(N_99), .Y(\data_from_adc[2]_69 ));
    CFG4 #( .INIT(16'h4000) )  \state_5_0_i_a2[1]  (.A(
        \state[0]_net_1 ), .B(N_54), .C(\cnt[5]_net_1 ), .D(
        \cnt[4]_net_1 ), .Y(N_86));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_8 (.A(freq_1), .B(
        \cnt_freq[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_7_net_1), .S(), .Y(), .FCO(cnt_freq6_cry_8_net_1)
        );
    SLE \freq[13]  (.D(freq15_net_1), .CLK(temp_sck_c), .EN(N_575_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(freq_6));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[6]  (.A(VCC_net_1), .B(
        \fpga_count[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[5]_net_1 ), .S(\fpga_count_s[6] ), .Y(), .FCO(
        \fpga_count_cry[6]_net_1 ));
    CFG4 #( .INIT(16'h5450) )  \temp_state_7_2_0_.N_11_i  (.A(m10_0_0), 
        .B(temp_count6), .C(\temp_state[0]_net_1 ), .D(
        \temp_state[1]_net_1 ), .Y(N_11_i_0));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_24 (.A(VCC_net_1), .B(
        temp_count[24]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_23_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_24_net_1));
    SLE \dac_count[2]  (.D(\dac_count_s[2] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[2]_net_1 ));
    SLE \cnt_freq[30]  (.D(\cnt_freq_s[30] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[30]_net_1 ));
    SLE \cnt_freq[29]  (.D(\cnt_freq_s[29] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[29]_net_1 ));
    SLE \fpga_shift_2[11]  (.D(BW_out_c[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[11]_net_1 ));
    SLE \fpga_data_receive[2]  (.D(BW_c[2]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[2]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNICB9I61[18]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[18]), .D(GND_net_1), .FCI(\temp_count_cry[17] ), .S(
        \temp_count_s[18] ), .Y(), .FCO(\temp_count_cry[18] ));
    SLE \cnt_freq[0]  (.D(\cnt_freq_s[0] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \cnt_frame_RNO_0[3]  (.A(cnt_frame_0_sqmuxa)
        , .Y(N_333_i));
    SLE \temp_count[24]  (.D(\temp_count_s[24] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[24]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9QGHR[12]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[12]), .D(GND_net_1), .FCI(\temp_count_cry[11] ), .S(
        \temp_count_s[12] ), .Y(), .FCO(\temp_count_cry[12] ));
    CFG4 #( .INIT(16'h1000) )  temp3_57_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_180), .Y(temp3_57));
    SLE \fpga_count[12]  (.D(\fpga_count_s[12] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[12]_net_1 ));
    CFG4 #( .INIT(16'hFEFA) )  \state_5_0_i_o4[1]  (.A(\cnt[3]_net_1 ), 
        .B(\cnt[1]_net_1 ), .C(\cnt[2]_net_1 ), .D(GPIO7_c), .Y(N_54));
    SLE \temp3[8]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_51), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[8]));
    CFG4 #( .INIT(16'h0080) )  \data_from_adc[2]_RNO_0[5]  (.A(GPIO7_c)
        , .B(\data_from_adc[2]_66_0_0_a2_0_out ), .C(\cnt[1]_net_1 ), 
        .D(\cnt[2]_net_1 ), .Y(\data_from_adc[2]_64_0_0_a2_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[6]  (.A(VCC_net_1), .B(
        \dac_count[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[5]_net_1 ), .S(\dac_count_s[6] ), .Y(), .FCO(
        \dac_count_cry[6]_net_1 ));
    SLE \temp2[2]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_29), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[2]));
    SLE \dac1_db[8]  (.D(N_705_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[8]));
    SLE \fpga_data_receive[14]  (.D(BW_c[14]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[14]_net_1 ));
    CFG3 #( .INIT(8'h12) )  \temp_count_data_RNO[1]  (.A(
        temp_count_data[0]), .B(temp_count_data[4]), .C(
        temp_count_data[1]), .Y(N_15_i_0));
    SLE \temp_count_data[1]  (.D(N_15_i_0), .CLK(temp_sck_c), .EN(
        N_17_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count_data[1]));
    SLE \state[1]  (.D(N_23_i_0), .CLK(temp_sck_c_i_0), .EN(N_70_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_15 (.A(freq_0), .B(
        \cnt_freq[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_14_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_15_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[13]  (.A(VCC_net_1), .B(
        \cnt_freq[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[12]_net_1 ), .S(\cnt_freq_s[13] ), .Y(), .FCO(
        \cnt_freq_cry[13]_net_1 ));
    CFG2 #( .INIT(4'h4) )  state15_0_a2 (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(state15));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9HN2C1[21]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[21]), .D(GND_net_1), .FCI(\temp_count_cry[20] ), .S(
        \temp_count_s[21] ), .Y(), .FCO(\temp_count_cry[21] ));
    CFG4 #( .INIT(16'h0040) )  \temp_count_data_RNO[4]  (.A(
        temp_count_data[4]), .B(temp_count_data[3]), .C(
        temp_count_data[2]), .D(N_76), .Y(N_6_i_0));
    CFG4 #( .INIT(16'h0100) )  freq3lto11 (.A(
        \data_from_adc[2][9]_net_1 ), .B(\data_from_adc[2][11]_net_1 ), 
        .C(\data_from_adc[2][10]_net_1 ), .D(freq3lt11), .Y(freq3));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[9]  (.A(
        \data_from_adc[2]_68_0_0_a2_0_out ), .B(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .C(
        \data_from_adc[2]_68_0_0_a2_0 ), .D(N_99), .Y(
        \data_from_adc[2]_68 ));
    SLE \cnt_freq[18]  (.D(\cnt_freq_s[18] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[18]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  temp3_52_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_180), .Y(temp3_52));
    ARI1 #( .INIT(20'h48421) )  fpga_flag4_0_I_15 (.A(
        \fpga_shift_2[11]_net_1 ), .B(\fpga_data_receive[10]_net_1 ), 
        .C(\fpga_data_receive[11]_net_1 ), .D(\fpga_shift_2[10]_net_1 )
        , .FCI(\fpga_flag4_0_data_tmp[4] ), .S(), .Y(), .FCO(
        \fpga_flag4_0_data_tmp[5] ));
    SLE \cnt[2]  (.D(\cnt_s[2] ), .CLK(temp_sck_c_i_0), .EN(cnte), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\cnt[2]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_26 (.A(VCC_net_1), .B(
        temp_count[26]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_25_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_26_net_1));
    SLE \data_from_adc[2][1]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_60 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][1]_net_1 ));
    ARI1 #( .INIT(20'h6AA00) )  cnt_freq6_cry_19 (.A(VCC_net_1), .B(
        \cnt_freq[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_18_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_19_net_1));
    ARI1 #( .INIT(20'h45500) )  temp_count6_cry_30 (.A(VCC_net_1), .B(
        temp_count[30]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_29_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_30_net_1));
    SLE \cnt_freq[14]  (.D(\cnt_freq_s[14] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[14]_net_1 ));
    CFG2 #( .INIT(4'h4) )  temp1_16_0_0_a2 (.A(temp_count_data[0]), .B(
        temp_count_data[1]), .Y(N_183));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[20]  (.A(VCC_net_1), .B(
        \cnt_freq[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[19]_net_1 ), .S(\cnt_freq_s[20] ), .Y(), .FCO(
        \cnt_freq_cry[20]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[29]  (.A(VCC_net_1), .B(
        \cnt_freq[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[28]_net_1 ), .S(\cnt_freq_s[29] ), .Y(), .FCO(
        \cnt_freq_cry[29]_net_1 ));
    SLE \temp3[0]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_43), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[0]));
    CFG4 #( .INIT(16'hFFF7) )  freq3lto8 (.A(
        \data_from_adc[2][7]_net_1 ), .B(\data_from_adc[2][8]_net_1 ), 
        .C(freq3lto8_1_net_1), .D(freq3lt8), .Y(freq3lt11));
    SLE \cnt_freq[12]  (.D(\cnt_freq_s[12] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[12]_net_1 ));
    SLE \temp1[12]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_23), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[12]));
    SLE \freq[16]  (.D(freq3), .CLK(temp_sck_c), .EN(N_575_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(freq_1));
    CFG4 #( .INIT(16'h0020) )  temp2_35_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_181), .D(N_76), .Y(temp2_35));
    SLE \dac_count[5]  (.D(\dac_count_s[5] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[5]_net_1 ));
    CFG4 #( .INIT(16'h1105) )  \state_RNO[0]  (.A(\state[0]_net_1 ), 
        .B(N_52), .C(GPIO11_c), .D(\state[1]_net_1 ), .Y(N_449_i_0));
    CFG1 #( .INIT(2'h1) )  \sdv_count_RNI847F[0]  (.A(
        \sdv_count[0]_net_1 ), .Y(\sdv_count_i_0[0] ));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[7]  (.A(VCC_net_1), .B(
        \dac_count[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[6]_net_1 ), .S(\dac_count_s[7] ), .Y(), .FCO(
        \dac_count_cry[7]_net_1 ));
    SLE \temp_count_data[3]  (.D(N_8_i_0), .CLK(temp_sck_c), .EN(
        N_17_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count_data[3]));
    CFG2 #( .INIT(4'h1) )  temp_count_data_n1_i_a2 (.A(
        temp_count_data[0]), .B(temp_count_data[1]), .Y(N_178));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_10 (.A(freq_0), .B(
        \cnt_freq[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_9_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_10_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_s[8]  (.A(VCC_net_1), .B(
        \dac_count[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[7]_net_1 ), .S(\dac_count_s[8]_net_1 ), .Y(), 
        .FCO());
    SLE GPIO14 (.D(fpga_flag_net_1), .CLK(BW_clk_c_i_0), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(GPIO14_c));
    SLE \cnt_freq[8]  (.D(\cnt_freq_s[8] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[8]_net_1 ));
    SLE \fpga_shift[8]  (.D(\fpga_count[8]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[8]));
    CFG1 #( .INIT(2'h1) )  \fpga_count_RNO[0]  (.A(
        \fpga_count[0]_net_1 ), .Y(\fpga_count_s[0] ));
    CFG4 #( .INIT(16'h6996) )  GPIO5_10 (.A(GPS2_Q0_c), .B(GPS2_LD_c), 
        .C(GPS1_Q1_c), .D(GPS1_Q0_c), .Y(GPIO5_10_net_1));
    SLE \dac1_db[9]  (.D(N_698_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[9]));
    CFG2 #( .INIT(4'h4) )  \cnt_RNI0B3K[5]  (.A(\cnt[5]_net_1 ), .B(
        \cnt_frame[1]_net_1 ), .Y(\data_from_adc[2]_59_0_0_a2_0_0 ));
    CFG4 #( .INIT(16'h0001) )  \SENSE_DOUT_1_RNO_0[1]  (.A(
        \cnt[5]_net_1 ), .B(\cnt[3]_net_1 ), .C(N_109), .D(
        \cnt[4]_net_1 ), .Y(N_39_i_0));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI6H37V[14]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[14]), .D(GND_net_1), .FCI(\temp_count_cry[13] ), .S(
        \temp_count_s[14] ), .Y(), .FCO(\temp_count_cry[14] ));
    ARI1 #( .INIT(20'h5AA55) )  temp_count6_cry_12 (.A(freq_2), .B(
        temp_count[12]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_11_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_12_net_1));
    SLE \fpga_count[14]  (.D(\fpga_count_s[14]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_count[14]_net_1 ));
    CFG4 #( .INIT(16'h0020) )  temp3_51_0_0_a3 (.A(temp_count_data[2]), 
        .B(temp_count_data[3]), .C(N_180), .D(N_76), .Y(temp3_51));
    ARI1 #( .INIT(20'h4AA00) )  cnt_freq_s_461 (.A(VCC_net_1), .B(
        \cnt_freq[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(cnt_freq_s_461_FCO));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIGDAQH[7]  (.A(VCC_net_1)
        , .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(temp_count[7]), .D(
        GND_net_1), .FCI(\temp_count_cry[6] ), .S(\temp_count_s[7] ), 
        .Y(), .FCO(\temp_count_cry[7] ));
    SLE \temp_count[7]  (.D(\temp_count_s[7] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[7]));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[5]  (.A(VCC_net_1), .B(
        \dac_count[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[4]_net_1 ), .S(\dac_count_s[5] ), .Y(), .FCO(
        \dac_count_cry[5]_net_1 ));
    SLE \temp_count[6]  (.D(\temp_count_s[6] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[6]));
    CFG3 #( .INIT(8'h80) )  \data_from_adc[2]_RNO[2]  (.A(N_99), .B(
        \data_from_adc[2]_66_0_0_a2_0_0 ), .C(\data_from_adc[2]_61_1 ), 
        .Y(\data_from_adc[2]_61 ));
    SLE \data_from_adc[2][0]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_59 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][0]_net_1 ));
    SLE \temp3[10]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_53), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[10]));
    SLE \data_from_adc[2][11]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_70 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][11]_net_1 ));
    SLE \temp_count[30]  (.D(\temp_count_s[30] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[30]));
    ARI1 #( .INIT(20'h4AA00) )  \dac_count_cry[3]  (.A(VCC_net_1), .B(
        \dac_count[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \dac_count_cry[2]_net_1 ), .S(\dac_count_s[3] ), .Y(), .FCO(
        \dac_count_cry[3]_net_1 ));
    CFG2 #( .INIT(4'h9) )  GPIO16_RNO (.A(cnt_freq6), .B(GPIO16_c), .Y(
        N_12_i_0));
    SLE \fpga_data_receive[9]  (.D(BW_c[9]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[9]_net_1 ));
    SLE \temp_count[31]  (.D(\temp_count_s[31] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[31]));
    SLE \cnt_frame[1]  (.D(cnt_frame_0), .CLK(temp_sck_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_frame[1]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_18 (.A(freq_11), .B(
        \cnt_freq[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_17_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_18_net_1));
    CFG2 #( .INIT(4'h1) )  clk_dac14 (.A(\sdv_count[1]_net_1 ), .B(
        \sdv_count[0]_net_1 ), .Y(clk_dac14_net_1));
    SLE \dac1_db[11]  (.D(N_684_i), .CLK(BW_clk_c), .EN(
        \sdv_count_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(dac1_db_c[11]));
    CFG4 #( .INIT(16'h8000) )  \un1_data_from_adc[2]_2lto11_i_a2_7  (
        .A(\data_from_adc[2][8]_net_1 ), .B(
        \data_from_adc[2][7]_net_1 ), .C(\data_from_adc[2][3]_net_1 ), 
        .D(\data_from_adc[2][2]_net_1 ), .Y(
        \un1_data_from_adc[2]_2lto11_i_a2_7_net_1 ));
    CFG4 #( .INIT(16'hC488) )  temp3_csn_RNO_0 (.A(
        \temp_state[2]_net_1 ), .B(\temp_state[0]_net_1 ), .C(
        temp_count_data[4]), .D(\temp_state[1]_net_1 ), .Y(
        un1_temp_state_7_or));
    CFG4 #( .INIT(16'h8000) )  \un1_data_from_adc[2]_2lto11_i_a2_6  (
        .A(\data_from_adc[2][4]_net_1 ), .B(
        \data_from_adc[2][11]_net_1 ), .C(\data_from_adc[2][6]_net_1 ), 
        .D(\data_from_adc[2][5]_net_1 ), .Y(
        \un1_data_from_adc[2]_2lto11_i_a2_6_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \un1_data_from_adc[2]_2lto11_i_a2_5  (
        .A(\data_from_adc[2][0]_net_1 ), .B(
        \data_from_adc[2][1]_net_1 ), .C(\data_from_adc[2][10]_net_1 ), 
        .D(\data_from_adc[2][9]_net_1 ), .Y(
        \un1_data_from_adc[2]_2lto11_i_a2_5_net_1 ));
    SLE \temp2[7]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_34), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[7]));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[4]  (.A(
        \data_from_adc[2]_66_0_0_a2_0_out ), .B(
        \data_from_adc[2]_63_0_0_a2_0 ), .C(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .D(N_99), .Y(
        \data_from_adc[2]_63 ));
    CFG2 #( .INIT(4'h7) )  \cnt_frame_0_0_o2[3]  (.A(
        \cnt_frame[0]_net_1 ), .B(\cnt_frame[1]_net_1 ), .Y(N_58));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[9]  (.A(VCC_net_1), .B(
        \fpga_count[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[8]_net_1 ), .S(\fpga_count_s[9] ), .Y(), .FCO(
        \fpga_count_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \fpga_count_cry[2]  (.A(VCC_net_1), .B(
        \fpga_count[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \fpga_count_cry[1]_net_1 ), .S(\fpga_count_s[2] ), .Y(), .FCO(
        \fpga_count_cry[2]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  temp1_13_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_182), .D(N_179), .Y(temp1_13));
    CFG4 #( .INIT(16'h8000) )  \data_from_adc[2]_RNO[3]  (.A(
        \data_from_adc[2]_70_0_0_a2_0 ), .B(N_99), .C(
        \data_from_adc[2]_66_0_0_a2_0_out ), .D(
        \data_from_adc[2]_59_0_0_a2_0_0 ), .Y(\data_from_adc[2]_62 ));
    SLE \temp2[10]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_37), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[10]));
    SLE \temp3[11]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp3_54), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp3[11]));
    SLE \temp_count[26]  (.D(\temp_count_s[26] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[26]));
    SLE \data_from_adc[2][7]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_66 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][7]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  temp2_40_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_181), .Y(temp2_40));
    SLE \fpga_shift_2[7]  (.D(BW_out_c[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[7]_net_1 ));
    SLE \data_from_adc[2][2]  (.D(GPIO4_c), .CLK(temp_sck_c), .EN(
        \data_from_adc[2]_61 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_from_adc[2][2]_net_1 ));
    SLE \dac_count[6]  (.D(\dac_count_s[6] ), .CLK(BW_clk_c), .EN(
        clk_dac14_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \dac_count[6]_net_1 ));
    SLE \cnt_freq[25]  (.D(\cnt_freq_s[25] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[25]_net_1 ));
    SLE \temp_count[18]  (.D(\temp_count_s[18] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[18]));
    SLE \temp1[7]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_18), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[7]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNILDBPQ1[29]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[29]), .D(GND_net_1), .FCI(\temp_count_cry[28] ), .S(
        \temp_count_s[29] ), .Y(), .FCO(\temp_count_cry[29] ));
    SLE temp2_csn (.D(temp2_csn_1_sqmuxa), .CLK(temp_sck_c), .EN(
        temp2_csn_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_322_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(temp2_csn_c));
    SLE \sdv_count[0]  (.D(\sdv_count_i_0[0] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\sdv_count[0]_net_1 ));
    CFG4 #( .INIT(16'h3500) )  \SENSE_DOUT_2_1_u_i_a2[1]  (.A(
        \cnt_frame[2]_net_1 ), .B(\cnt[1]_net_1 ), .C(\cnt[2]_net_1 ), 
        .D(\SENSE_DOUT_2_1_u_i_a2_0[1]_net_1 ), .Y(N_80));
    CFG3 #( .INIT(8'h08) )  \cnt_RNIBCML_1[1]  (.A(\cnt[2]_net_1 ), .B(
        GPIO7_c), .C(\cnt[1]_net_1 ), .Y(
        \data_from_adc[2]_70_0_0_a2_0 ));
    SLE \temp_count[3]  (.D(\temp_count_s[3] ), .CLK(temp_sck_c), .EN(
        \temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(temp_count[3]));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNI9NR8L1[26]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[26]), .D(GND_net_1), .FCI(\temp_count_cry[25] ), .S(
        \temp_count_s[26] ), .Y(), .FCO(\temp_count_cry[26] ));
    SLE \fpga_shift[5]  (.D(\fpga_count[5]_net_1 ), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(BW_out_c[5]));
    SLE \fpga_count[0]  (.D(\fpga_count_s[0] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[0]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \temp_count_RNIGQGUO1[28]  (.A(
        VCC_net_1), .B(temp_count6_cry_31_RNIPJ5K1_Y), .C(
        temp_count[28]), .D(GND_net_1), .FCI(\temp_count_cry[27] ), .S(
        \temp_count_s[28] ), .Y(), .FCO(\temp_count_cry[28] ));
    ARI1 #( .INIT(20'h6AA00) )  temp_count6_cry_19 (.A(VCC_net_1), .B(
        temp_count[19]), .C(GND_net_1), .D(GND_net_1), .FCI(
        temp_count6_cry_18_net_1), .S(), .Y(), .FCO(
        temp_count6_cry_19_net_1));
    SLE \freq[21]  (.D(N_445_i_0), .CLK(temp_sck_c), .EN(N_575_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(freq_14));
    SLE \fpga_count[4]  (.D(\fpga_count_s[4] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[4]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  temp1_20_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_179), .Y(temp1_20));
    CFG4 #( .INIT(16'h2000) )  temp1_16_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_179), .Y(temp1_16));
    SLE \temp1[14]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_25), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[14]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[18]  (.A(VCC_net_1), .B(
        \cnt_freq[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[17]_net_1 ), .S(\cnt_freq_s[18] ), .Y(), .FCO(
        \cnt_freq_cry[18]_net_1 ));
    SLE \cnt_freq[20]  (.D(\cnt_freq_s[20] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[20]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[16]  (.A(VCC_net_1), .B(
        \cnt_freq[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[15]_net_1 ), .S(\cnt_freq_s[16] ), .Y(), .FCO(
        \cnt_freq_cry[16]_net_1 ));
    SLE \temp2[11]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp2_38), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp2[11]));
    ARI1 #( .INIT(20'h4AA00) )  \cnt_freq_cry[5]  (.A(VCC_net_1), .B(
        \cnt_freq[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \cnt_freq_cry[4]_net_1 ), .S(\cnt_freq_s[5] ), .Y(), .FCO(
        \cnt_freq_cry[5]_net_1 ));
    SLE \cnt_freq[27]  (.D(\cnt_freq_s[27] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[27]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  temp3_48_0_0_a3 (.A(temp_count_data[3]), 
        .B(temp_count_data[2]), .C(N_183), .D(N_180), .Y(temp3_48));
    CFG2 #( .INIT(4'hE) )  temp1_csn_RNO (.A(temp_state26), .B(
        un1_temp_state_8_or), .Y(temp1_csn_RNO_net_1));
    CFG4 #( .INIT(16'h6996) )  GPIO3 (.A(GPIO3_9_net_1), .B(
        GPIO3_8_net_1), .C(GPIO3_7_net_1), .D(GPIO3_6_net_1), .Y(
        GPIO3_c));
    CFG4 #( .INIT(16'h0400) )  \cnt_frame_0_0_a2_0_2[3]  (.A(
        \state[1]_net_1 ), .B(\cnt_frame[2]_net_1 ), .C(N_58), .D(
        \state[0]_net_1 ), .Y(\cnt_frame_0_0_a2_0_2[3]_net_1 ));
    SLE SENSE_CS_1 (.D(N_21), .CLK(temp_sck_c_i_0), .EN(state15), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(SENSE_CS_1_c));
    SLE \fpga_data_receive[7]  (.D(BW_c[7]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[7]_net_1 ));
    CFG4 #( .INIT(16'h3222) )  clk_dac1_2 (.A(\sdv_count_i_0[1] ), .B(
        clk_dac14_net_1), .C(dac1_clk_c), .D(\sdv_count[1]_net_1 ), .Y(
        clk_dac1_2_net_1));
    SLE \fpga_count[11]  (.D(\fpga_count_s[11] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_count[11]_net_1 ));
    SLE \temp1[3]  (.D(temp_so_c), .CLK(temp_sck_c), .EN(temp1_14), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(temp1[3]));
    SLE \fpga_shift_2[10]  (.D(BW_out_c[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fpga_shift_2[10]_net_1 ));
    SLE \fpga_data_receive[4]  (.D(BW_c[4]), .CLK(BW_clk_c_i_0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fpga_data_receive[4]_net_1 ));
    CFG2 #( .INIT(4'hE) )  temp2_csn_RNO (.A(temp_state26), .B(
        un1_temp_state29_3_or), .Y(temp2_csn_RNO_net_1));
    SLE \cnt_freq[1]  (.D(\cnt_freq_s[1] ), .CLK(temp_sck_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(cnt_freq6), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\cnt_freq[1]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_13 (.A(freq_6), .B(
        \cnt_freq[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_12_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_13_net_1));
    ARI1 #( .INIT(20'h5AA55) )  cnt_freq6_cry_11 (.A(freq_1), .B(
        \cnt_freq[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        cnt_freq6_cry_10_net_1), .S(), .Y(), .FCO(
        cnt_freq6_cry_11_net_1));
    CFG2 #( .INIT(4'h1) )  temp_count_data_n0_i_a3 (.A(
        temp_count_data[4]), .B(temp_count_data[0]), .Y(N_113));
    SLE \temp_count[23]  (.D(\temp_count_s[23] ), .CLK(temp_sck_c), 
        .EN(\temp_state_i_0[0] ), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        temp_count[23]));
    
endmodule


module b5_nvmFL_465s_x_0(
       b4_nUAi,
       IICE_comm2iice,
       b4_PLyF,
       b7_PSyi3wy,
       b8_PSyiBgYG
    );
output [463:0] b4_nUAi;
input  [11:10] IICE_comm2iice;
input  b4_PLyF;
output b7_PSyi3wy;
input  b8_PSyiBgYG;

    wire VCC_net_1, b6_OKctIF4_net_1, GND_net_1;
    
    SLE \b6_OKctIF[169]  (.D(b4_nUAi[294]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[295]));
    SLE \b6_OKctIF[41]  (.D(b4_nUAi[422]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[423]));
    SLE \b6_OKctIF[269]  (.D(b4_nUAi[194]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[195]));
    SLE \b6_OKctIF[147]  (.D(b4_nUAi[316]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[317]));
    SLE \b6_OKctIF[58]  (.D(b4_nUAi[405]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[406]));
    SLE \b6_OKctIF[55]  (.D(b4_nUAi[408]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[409]));
    SLE \b6_OKctIF[352]  (.D(b4_nUAi[111]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[112]));
    SLE \b6_OKctIF[430]  (.D(b4_nUAi[33]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[34]));
    SLE \b6_OKctIF[204]  (.D(b4_nUAi[259]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[260]));
    SLE \b6_OKctIF[374]  (.D(b4_nUAi[89]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[90]));
    SLE \b6_OKctIF[284]  (.D(b4_nUAi[179]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[180]));
    SLE \b6_OKctIF[2]  (.D(b4_nUAi[461]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[462]));
    SLE \b6_OKctIF[260]  (.D(b4_nUAi[203]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[204]));
    SLE \b6_OKctIF[156]  (.D(b4_nUAi[307]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[308]));
    SLE \b6_OKctIF[47]  (.D(b4_nUAi[416]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[417]));
    SLE \b6_OKctIF[212]  (.D(b4_nUAi[251]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[252]));
    SLE \b6_OKctIF[165]  (.D(b4_nUAi[298]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[299]));
    SLE \b6_OKctIF[46]  (.D(b4_nUAi[417]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[418]));
    SLE \b6_OKctIF[43]  (.D(b4_nUAi[420]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[421]));
    SLE \b6_OKctIF[208]  (.D(b4_nUAi[255]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[256]));
    SLE \b6_OKctIF[288]  (.D(b4_nUAi[175]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[176]));
    SLE \b6_OKctIF[405]  (.D(b4_nUAi[58]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[59]));
    SLE \b6_OKctIF[246]  (.D(b4_nUAi[217]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[218]));
    SLE \b6_OKctIF[312]  (.D(b4_nUAi[151]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[152]));
    SLE \b6_OKctIF[251]  (.D(b4_nUAi[212]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[213]));
    SLE \b6_OKctIF[116]  (.D(b4_nUAi[347]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[348]));
    SLE \b6_OKctIF[409]  (.D(b4_nUAi[54]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[55]));
    CFG2 #( .INIT(4'h8) )  b6_OKctIF4 (.A(b8_PSyiBgYG), .B(
        IICE_comm2iice[10]), .Y(b6_OKctIF4_net_1));
    SLE \b6_OKctIF[401]  (.D(b4_nUAi[62]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[63]));
    SLE \b6_OKctIF[334]  (.D(b4_nUAi[129]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[130]));
    SLE \b6_OKctIF[428]  (.D(b4_nUAi[35]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[36]));
    SLE \b6_OKctIF[341]  (.D(b4_nUAi[122]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[123]));
    SLE \b6_OKctIF[211]  (.D(b4_nUAi[252]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[253]));
    SLE \b6_OKctIF[100]  (.D(b4_nUAi[363]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[364]));
    SLE \b6_OKctIF[437]  (.D(b4_nUAi[26]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[27]));
    SLE \b6_OKctIF[42]  (.D(b4_nUAi[421]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[422]));
    SLE \b6_OKctIF[348]  (.D(b4_nUAi[115]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[116]));
    SLE \b6_OKctIF[194]  (.D(b4_nUAi[269]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[270]));
    SLE \b6_OKctIF[180]  (.D(b4_nUAi[283]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[284]));
    SLE \b6_OKctIF[403]  (.D(b4_nUAi[60]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[61]));
    SLE \b6_OKctIF[432]  (.D(b4_nUAi[31]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[32]));
    SLE \b6_OKctIF[375]  (.D(b4_nUAi[88]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[89]));
    SLE \b6_OKctIF[275]  (.D(b4_nUAi[188]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[189]));
    SLE \b6_OKctIF[49]  (.D(b4_nUAi[414]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[415]));
    SLE \b6_OKctIF[377]  (.D(b4_nUAi[86]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[87]));
    SLE \b6_OKctIF[390]  (.D(b4_nUAi[73]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[74]));
    SLE \b6_OKctIF[103]  (.D(b4_nUAi[360]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[361]));
    SLE \b6_OKctIF[183]  (.D(b4_nUAi[280]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[281]));
    SLE \b6_OKctIF[440]  (.D(b4_nUAi[23]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[24]));
    SLE \b6_OKctIF[124]  (.D(b4_nUAi[339]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[340]));
    SLE \b6_OKctIF[264]  (.D(b4_nUAi[199]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[200]));
    SLE \b6_OKctIF[197]  (.D(b4_nUAi[266]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[267]));
    SLE \b6_OKctIF[102]  (.D(b4_nUAi[361]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[362]));
    SLE \b6_OKctIF[320]  (.D(b4_nUAi[143]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[144]));
    SLE \b6_OKctIF[182]  (.D(b4_nUAi[281]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[282]));
    SLE \b6_OKctIF[40]  (.D(b4_nUAi[423]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[424]));
    SLE \b6_OKctIF[268]  (.D(b4_nUAi[195]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[196]));
    SLE \b6_OKctIF[127]  (.D(b4_nUAi[336]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[337]));
    SLE \b6_OKctIF[458]  (.D(b4_nUAi[5]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[6]));
    SLE \b6_OKctIF[3]  (.D(b4_nUAi[460]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[461]));
    SLE \b6_OKctIF[296]  (.D(b4_nUAi[167]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[168]));
    SLE \b6_OKctIF[335]  (.D(b4_nUAi[128]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[129]));
    SLE \b6_OKctIF[235]  (.D(b4_nUAi[228]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[229]));
    SLE \b6_OKctIF[337]  (.D(b4_nUAi[126]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[127]));
    SLE \b6_OKctIF[154]  (.D(b4_nUAi[309]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[310]));
    SLE \b6_OKctIF[226]  (.D(b4_nUAi[237]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[238]));
    SLE \b6_OKctIF[461]  (.D(b4_nUAi[2]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[3]));
    SLE \b6_OKctIF[418]  (.D(b4_nUAi[45]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[46]));
    SLE \b6_OKctIF[344]  (.D(b4_nUAi[119]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[120]));
    SLE \b6_OKctIF[350]  (.D(b4_nUAi[113]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[114]));
    SLE \b6_OKctIF[447]  (.D(b4_nUAi[16]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[17]));
    SLE \b6_OKctIF[160]  (.D(b4_nUAi[303]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[304]));
    SLE \b6_OKctIF[404]  (.D(b4_nUAi[59]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[60]));
    SLE \b6_OKctIF[24]  (.D(b4_nUAi[439]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[440]));
    SLE \b6_OKctIF[463]  (.D(b4_nUAi[0]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[1]));
    SLE \b6_OKctIF[442]  (.D(b4_nUAi[21]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[22]));
    SLE \b6_OKctIF[178]  (.D(b4_nUAi[285]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[286]));
    SLE \b6_OKctIF[391]  (.D(b4_nUAi[72]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[73]));
    SLE \b6_OKctIF[157]  (.D(b4_nUAi[306]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[307]));
    SLE \b6_OKctIF[398]  (.D(b4_nUAi[65]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[66]));
    SLE \b6_OKctIF[163]  (.D(b4_nUAi[300]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[301]));
    SLE \b6_OKctIF[114]  (.D(b4_nUAi[349]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[350]));
    GND GND (.Y(GND_net_1));
    SLE \b6_OKctIF[21]  (.D(b4_nUAi[442]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[443]));
    SLE \b6_OKctIF[321]  (.D(b4_nUAi[142]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[143]));
    SLE \b6_OKctIF[310]  (.D(b4_nUAi[153]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[154]));
    SLE \b6_OKctIF[328]  (.D(b4_nUAi[135]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[136]));
    SLE \b6_OKctIF[162]  (.D(b4_nUAi[301]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[302]));
    SLE \b6_OKctIF[5]  (.D(b4_nUAi[458]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[459]));
    SLE \b6_OKctIF[27]  (.D(b4_nUAi[436]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[437]));
    SLE \b6_OKctIF[207]  (.D(b4_nUAi[256]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[257]));
    SLE \b6_OKctIF[287]  (.D(b4_nUAi[176]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[177]));
    SLE \b6_OKctIF[256]  (.D(b4_nUAi[207]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[208]));
    SLE \b6_OKctIF[54]  (.D(b4_nUAi[409]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[410]));
    SLE \b6_OKctIF[273]  (.D(b4_nUAi[190]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[191]));
    SLE \b6_OKctIF[117]  (.D(b4_nUAi[346]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[347]));
    SLE \b6_OKctIF[26]  (.D(b4_nUAi[437]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[438]));
    SLE \b6_OKctIF[23]  (.D(b4_nUAi[440]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[441]));
    SLE \b6_OKctIF[373]  (.D(b4_nUAi[90]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[91]));
    SLE \b6_OKctIF[420]  (.D(b4_nUAi[43]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[44]));
    SLE \b6_OKctIF[376]  (.D(b4_nUAi[87]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[88]));
    SLE \b6_OKctIF[171]  (.D(b4_nUAi[292]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[293]));
    SLE \b6_OKctIF[51]  (.D(b4_nUAi[412]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[413]));
    SLE \b6_OKctIF[345]  (.D(b4_nUAi[118]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[119]));
    SLE \b6_OKctIF[245]  (.D(b4_nUAi[218]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[219]));
    SLE \b6_OKctIF[138]  (.D(b4_nUAi[325]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[326]));
    SLE \b6_OKctIF[347]  (.D(b4_nUAi[116]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[117]));
    SLE \b6_OKctIF[216]  (.D(b4_nUAi[247]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[248]));
    SLE \b6_OKctIF[57]  (.D(b4_nUAi[406]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[407]));
    SLE \b6_OKctIF[351]  (.D(b4_nUAi[112]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[113]));
    SLE \b6_OKctIF[56]  (.D(b4_nUAi[407]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[408]));
    SLE \b6_OKctIF[53]  (.D(b4_nUAi[410]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[411]));
    SLE \b6_OKctIF[358]  (.D(b4_nUAi[105]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[106]));
    SLE \b6_OKctIF[202]  (.D(b4_nUAi[261]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[262]));
    SLE \b6_OKctIF[38]  (.D(b4_nUAi[425]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[426]));
    SLE \b6_OKctIF[35]  (.D(b4_nUAi[428]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[429]));
    SLE \b6_OKctIF[282]  (.D(b4_nUAi[181]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[182]));
    SLE \b6_OKctIF[464]  (.D(b4_PLyF), .CLK(IICE_comm2iice[11]), .EN(
        b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[0]));
    SLE \b6_OKctIF[394]  (.D(b4_nUAi[69]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[70]));
    SLE \b6_OKctIF[22]  (.D(b4_nUAi[441]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[442]));
    SLE \b6_OKctIF[233]  (.D(b4_nUAi[230]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[231]));
    SLE \b6_OKctIF[333]  (.D(b4_nUAi[130]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[131]));
    SLE \b6_OKctIF[29]  (.D(b4_nUAi[434]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[435]));
    SLE \b6_OKctIF[450]  (.D(b4_nUAi[13]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[14]));
    SLE \b6_OKctIF[302]  (.D(b4_nUAi[161]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[162]));
    SLE \b6_OKctIF[382]  (.D(b4_nUAi[81]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[82]));
    SLE \b6_OKctIF[336]  (.D(b4_nUAi[127]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[128]));
    SLE \b6_OKctIF[324]  (.D(b4_nUAi[139]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[140]));
    SLE \b6_OKctIF[311]  (.D(b4_nUAi[152]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[153]));
    SLE \b6_OKctIF[131]  (.D(b4_nUAi[332]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[333]));
    SLE \b6_OKctIF[106]  (.D(b4_nUAi[357]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[358]));
    SLE \b6_OKctIF[9]  (.D(b4_nUAi[454]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[455]));
    SLE \b6_OKctIF[318]  (.D(b4_nUAi[145]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[146]));
    SLE \b6_OKctIF[186]  (.D(b4_nUAi[277]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[278]));
    SLE \b6_OKctIF[427]  (.D(b4_nUAi[36]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[37]));
    SLE \b6_OKctIF[422]  (.D(b4_nUAi[41]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[42]));
    SLE \b6_OKctIF[379]  (.D(b4_nUAi[84]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[85]));
    SLE \b6_OKctIF[267]  (.D(b4_nUAi[196]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[197]));
    SLE \b6_OKctIF[20]  (.D(b4_nUAi[443]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[444]));
    SLE \b6_OKctIF[52]  (.D(b4_nUAi[411]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[412]));
    SLE \b6_OKctIF[410]  (.D(b4_nUAi[53]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[54]));
    SLE \b6_OKctIF[201]  (.D(b4_nUAi[262]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[263]));
    SLE \b6_OKctIF[179]  (.D(b4_nUAi[284]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[285]));
    SLE \b6_OKctIF[59]  (.D(b4_nUAi[404]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[405]));
    SLE \b6_OKctIF[281]  (.D(b4_nUAi[182]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[183]));
    SLE \b6_OKctIF[279]  (.D(b4_nUAi[184]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[185]));
    SLE \b6_OKctIF[148]  (.D(b4_nUAi[315]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[316]));
    SLE \b6_OKctIF[18]  (.D(b4_nUAi[445]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[446]));
    SLE \b6_OKctIF[15]  (.D(b4_nUAi[448]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[449]));
    SLE \b6_OKctIF[270]  (.D(b4_nUAi[193]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[194]));
    SLE \b6_OKctIF[395]  (.D(b4_nUAi[68]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[69]));
    SLE \b6_OKctIF[295]  (.D(b4_nUAi[168]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[169]));
    SLE \b6_OKctIF[175]  (.D(b4_nUAi[288]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[289]));
    SLE \b6_OKctIF[397]  (.D(b4_nUAi[66]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[67]));
    SLE \b6_OKctIF[354]  (.D(b4_nUAi[109]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[110]));
    VCC VCC (.Y(VCC_net_1));
    SLE \b6_OKctIF[50]  (.D(b4_nUAi[413]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[414]));
    SLE \b6_OKctIF[457]  (.D(b4_nUAi[6]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[7]));
    SLE \b6_OKctIF[262]  (.D(b4_nUAi[201]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[202]));
    SLE \b6_OKctIF[452]  (.D(b4_nUAi[11]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[12]));
    SLE \b6_OKctIF[78]  (.D(b4_nUAi[385]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[386]));
    SLE \b6_OKctIF[75]  (.D(b4_nUAi[388]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[389]));
    SLE \b6_OKctIF[339]  (.D(b4_nUAi[124]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[125]));
    SLE \b6_OKctIF[325]  (.D(b4_nUAi[138]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[139]));
    SLE \b6_OKctIF[225]  (.D(b4_nUAi[238]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[239]));
    SLE \b6_OKctIF[327]  (.D(b4_nUAi[136]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[137]));
    SLE \b6_OKctIF[436]  (.D(b4_nUAi[27]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[28]));
    SLE \b6_OKctIF[243]  (.D(b4_nUAi[220]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[221]));
    SLE \b6_OKctIF[343]  (.D(b4_nUAi[120]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[121]));
    SLE \b6_OKctIF[68]  (.D(b4_nUAi[395]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[396]));
    SLE \b6_OKctIF[65]  (.D(b4_nUAi[398]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[399]));
    SLE \b6_OKctIF[362]  (.D(b4_nUAi[101]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[102]));
    SLE \b6_OKctIF[139]  (.D(b4_nUAi[324]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[325]));
    SLE \b6_OKctIF[314]  (.D(b4_nUAi[149]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[150]));
    SLE \b6_OKctIF[239]  (.D(b4_nUAi[224]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[225]));
    SLE \b6_OKctIF[346]  (.D(b4_nUAi[117]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[118]));
    SLE \b6_OKctIF[141]  (.D(b4_nUAi[322]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[323]));
    SLE \b6_OKctIF[417]  (.D(b4_nUAi[46]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[47]));
    SLE \b6_OKctIF[166]  (.D(b4_nUAi[297]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[298]));
    SLE \b6_OKctIF[412]  (.D(b4_nUAi[51]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[52]));
    SLE \b6_OKctIF[230]  (.D(b4_nUAi[233]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[234]));
    SLE \b6_OKctIF[135]  (.D(b4_nUAi[328]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[329]));
    SLE \b6_OKctIF[408]  (.D(b4_nUAi[55]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[56]));
    SLE \b6_OKctIF[261]  (.D(b4_nUAi[202]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[203]));
    SLE \b6_OKctIF[355]  (.D(b4_nUAi[108]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[109]));
    SLE \b6_OKctIF[255]  (.D(b4_nUAi[208]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[209]));
    SLE \b6_OKctIF[357]  (.D(b4_nUAi[106]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[107]));
    SLE \b6_OKctIF[98]  (.D(b4_nUAi[365]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[366]));
    SLE \b6_OKctIF[95]  (.D(b4_nUAi[368]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[369]));
    SLE \b6_OKctIF[274]  (.D(b4_nUAi[189]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[190]));
    SLE \b6_OKctIF[198]  (.D(b4_nUAi[265]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[266]));
    SLE \b6_OKctIF[104]  (.D(b4_nUAi[359]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[360]));
    SLE \b6_OKctIF[184]  (.D(b4_nUAi[279]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[280]));
    SLE \b6_OKctIF[278]  (.D(b4_nUAi[185]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[186]));
    SLE \b6_OKctIF[300]  (.D(b4_nUAi[163]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[164]));
    SLE \b6_OKctIF[380]  (.D(b4_nUAi[83]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[84]));
    SLE \b6_OKctIF[315]  (.D(b4_nUAi[148]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[149]));
    SLE \b6_OKctIF[215]  (.D(b4_nUAi[248]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[249]));
    SLE \b6_OKctIF[349]  (.D(b4_nUAi[114]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[115]));
    SLE \b6_OKctIF[317]  (.D(b4_nUAi[146]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[147]));
    SLE \b6_OKctIF[128]  (.D(b4_nUAi[335]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[336]));
    SLE \b6_OKctIF[446]  (.D(b4_nUAi[17]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[18]));
    SLE \b6_OKctIF[107]  (.D(b4_nUAi[356]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[357]));
    SLE \b6_OKctIF[187]  (.D(b4_nUAi[276]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[277]));
    SLE \b6_OKctIF[149]  (.D(b4_nUAi[314]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[315]));
    SLE \b6_OKctIF[293]  (.D(b4_nUAi[170]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[171]));
    SLE \b6_OKctIF[249]  (.D(b4_nUAi[214]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[215]));
    SLE \b6_OKctIF[393]  (.D(b4_nUAi[70]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[71]));
    SLE \b6_OKctIF[34]  (.D(b4_nUAi[429]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[430]));
    SLE \b6_OKctIF[7]  (.D(b4_nUAi[456]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[457]));
    SLE \b6_OKctIF[234]  (.D(b4_nUAi[229]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[230]));
    SLE \b6_OKctIF[396]  (.D(b4_nUAi[67]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[68]));
    SLE \b6_OKctIF[240]  (.D(b4_nUAi[223]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[224]));
    SLE \b6_OKctIF[191]  (.D(b4_nUAi[272]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[273]));
    SLE \b6_OKctIF[206]  (.D(b4_nUAi[257]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[258]));
    SLE \b6_OKctIF[145]  (.D(b4_nUAi[318]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[319]));
    SLE \b6_OKctIF[286]  (.D(b4_nUAi[177]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[178]));
    SLE \b6_OKctIF[223]  (.D(b4_nUAi[240]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[241]));
    SLE \b6_OKctIF[170]  (.D(b4_nUAi[293]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[294]));
    SLE \b6_OKctIF[88]  (.D(b4_nUAi[375]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[376]));
    SLE \b6_OKctIF[85]  (.D(b4_nUAi[378]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[379]));
    SLE \b6_OKctIF[6]  (.D(b4_nUAi[457]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[458]));
    SLE \b6_OKctIF[31]  (.D(b4_nUAi[432]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[433]));
    SLE \b6_OKctIF[323]  (.D(b4_nUAi[140]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[141]));
    SLE \b6_OKctIF[238]  (.D(b4_nUAi[225]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[226]));
    SLE \b6_OKctIF[435]  (.D(b4_nUAi[28]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[29]));
    SLE \b6_OKctIF[326]  (.D(b4_nUAi[137]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[138]));
    SLE \b6_OKctIF[173]  (.D(b4_nUAi[290]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[291]));
    SLE \b6_OKctIF[158]  (.D(b4_nUAi[305]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[306]));
    SLE \b6_OKctIF[121]  (.D(b4_nUAi[342]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[343]));
    SLE \b6_OKctIF[37]  (.D(b4_nUAi[426]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[427]));
    SLE \b6_OKctIF[36]  (.D(b4_nUAi[427]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[428]));
    SLE \b6_OKctIF[33]  (.D(b4_nUAi[430]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[431]));
    SLE \b6_OKctIF[172]  (.D(b4_nUAi[291]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[292]));
    SLE \b6_OKctIF[164]  (.D(b4_nUAi[299]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[300]));
    SLE \b6_OKctIF[439]  (.D(b4_nUAi[24]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[25]));
    SLE \b6_OKctIF[4]  (.D(b4_nUAi[459]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[460]));
    SLE \b6_OKctIF[301]  (.D(b4_nUAi[162]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[163]));
    SLE \b6_OKctIF[381]  (.D(b4_nUAi[82]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[83]));
    SLE \b6_OKctIF[308]  (.D(b4_nUAi[155]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[156]));
    SLE \b6_OKctIF[388]  (.D(b4_nUAi[75]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[76]));
    SLE \b6_OKctIF[360]  (.D(b4_nUAi[103]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[104]));
    SLE \b6_OKctIF[431]  (.D(b4_nUAi[32]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[33]));
    SLE \b6_OKctIF[118]  (.D(b4_nUAi[345]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[346]));
    SLE \b6_OKctIF[14]  (.D(b4_nUAi[449]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[450]));
    SLE \b6_OKctIF[253]  (.D(b4_nUAi[210]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[211]));
    SLE \b6_OKctIF[130]  (.D(b4_nUAi[333]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[334]));
    SLE \b6_OKctIF[353]  (.D(b4_nUAi[110]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[111]));
    SLE \b6_OKctIF[167]  (.D(b4_nUAi[296]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[297]));
    SLE \b6_OKctIF[433]  (.D(b4_nUAi[30]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[31]));
    SLE \b6_OKctIF[400]  (.D(b4_nUAi[63]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[64]));
    SLE \b6_OKctIF[399]  (.D(b4_nUAi[64]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[65]));
    SLE \b6_OKctIF[356]  (.D(b4_nUAi[107]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[108]));
    SLE \b6_OKctIF[151]  (.D(b4_nUAi[312]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[313]));
    SLE \b6_OKctIF[11]  (.D(b4_nUAi[452]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[453]));
    SLE \b6_OKctIF[133]  (.D(b4_nUAi[330]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[331]));
    SLE \b6_OKctIF[74]  (.D(b4_nUAi[389]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[390]));
    SLE \b6_OKctIF[32]  (.D(b4_nUAi[431]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[432]));
    SLE \b6_OKctIF[199]  (.D(b4_nUAi[264]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[265]));
    SLE \b6_OKctIF[299]  (.D(b4_nUAi[164]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[165]));
    SLE \b6_OKctIF[244]  (.D(b4_nUAi[219]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[220]));
    SLE \b6_OKctIF[329]  (.D(b4_nUAi[134]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[135]));
    SLE \b6_OKctIF[39]  (.D(b4_nUAi[424]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[425]));
    SLE \b6_OKctIF[213]  (.D(b4_nUAi[250]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[251]));
    SLE \b6_OKctIF[17]  (.D(b4_nUAi[446]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[447]));
    SLE \b6_OKctIF[426]  (.D(b4_nUAi[37]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[38]));
    SLE \b6_OKctIF[266]  (.D(b4_nUAi[197]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[198]));
    SLE \b6_OKctIF[132]  (.D(b4_nUAi[331]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[332]));
    SLE \b6_OKctIF[64]  (.D(b4_nUAi[399]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[400]));
    SLE \b6_OKctIF[313]  (.D(b4_nUAi[150]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[151]));
    SLE \b6_OKctIF[16]  (.D(b4_nUAi[447]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[448]));
    SLE \b6_OKctIF[13]  (.D(b4_nUAi[450]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[451]));
    SLE \b6_OKctIF[71]  (.D(b4_nUAi[392]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[393]));
    SLE \b6_OKctIF[290]  (.D(b4_nUAi[173]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[174]));
    SLE \b6_OKctIF[248]  (.D(b4_nUAi[215]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[216]));
    SLE \b6_OKctIF[195]  (.D(b4_nUAi[268]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[269]));
    SLE \b6_OKctIF[129]  (.D(b4_nUAi[334]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[335]));
    SLE \b6_OKctIF[445]  (.D(b4_nUAi[18]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[19]));
    SLE \b6_OKctIF[316]  (.D(b4_nUAi[147]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[148]));
    SLE \b6_OKctIF[229]  (.D(b4_nUAi[234]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[235]));
    SLE \b6_OKctIF[111]  (.D(b4_nUAi[352]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[353]));
    SLE \b6_OKctIF[61]  (.D(b4_nUAi[402]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[403]));
    SLE \b6_OKctIF[77]  (.D(b4_nUAi[386]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[387]));
    SLE \b6_OKctIF[30]  (.D(b4_nUAi[433]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[434]));
    SLE \b6_OKctIF[220]  (.D(b4_nUAi[243]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[244]));
    SLE \b6_OKctIF[125]  (.D(b4_nUAi[338]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[339]));
    SLE \b6_OKctIF[76]  (.D(b4_nUAi[387]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[388]));
    SLE \b6_OKctIF[73]  (.D(b4_nUAi[390]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[391]));
    SLE \b6_OKctIF[449]  (.D(b4_nUAi[14]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[15]));
    SLE \b6_OKctIF[304]  (.D(b4_nUAi[159]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[160]));
    SLE \b6_OKctIF[67]  (.D(b4_nUAi[396]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[397]));
    SLE \b6_OKctIF[384]  (.D(b4_nUAi[79]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[80]));
    SLE \b6_OKctIF[361]  (.D(b4_nUAi[102]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[103]));
    SLE \b6_OKctIF[277]  (.D(b4_nUAi[186]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[187]));
    SLE \b6_OKctIF[407]  (.D(b4_nUAi[56]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[57]));
    SLE \b6_OKctIF[66]  (.D(b4_nUAi[397]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[398]));
    SLE \b6_OKctIF[63]  (.D(b4_nUAi[400]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[401]));
    SLE \b6_OKctIF[368]  (.D(b4_nUAi[95]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[96]));
    SLE \b6_OKctIF[441]  (.D(b4_nUAi[22]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[23]));
    SLE \b6_OKctIF[402]  (.D(b4_nUAi[61]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[62]));
    SLE \b6_OKctIF[359]  (.D(b4_nUAi[104]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[105]));
    SLE \b6_OKctIF[94]  (.D(b4_nUAi[369]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[370]));
    SLE \b6_OKctIF[456]  (.D(b4_nUAi[7]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[8]));
    SLE \b6_OKctIF[140]  (.D(b4_nUAi[323]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[324]));
    SLE \b6_OKctIF[12]  (.D(b4_nUAi[451]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[452]));
    SLE \b6_OKctIF[443]  (.D(b4_nUAi[20]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[21]));
    SLE \b6_OKctIF[434]  (.D(b4_nUAi[29]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[30]));
    SLE \b6_OKctIF[19]  (.D(b4_nUAi[444]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[445]));
    SLE \b6_OKctIF[159]  (.D(b4_nUAi[304]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[305]));
    SLE \b6_OKctIF[460]  (.D(b4_nUAi[3]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[4]));
    SLE \b6_OKctIF[259]  (.D(b4_nUAi[204]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[205]));
    SLE \b6_OKctIF[91]  (.D(b4_nUAi[372]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[373]));
    SLE \b6_OKctIF[143]  (.D(b4_nUAi[320]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[321]));
    SLE \b6_OKctIF[319]  (.D(b4_nUAi[144]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[145]));
    SLE \b6_OKctIF[250]  (.D(b4_nUAi[213]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[214]));
    SLE \b6_OKctIF[72]  (.D(b4_nUAi[391]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[392]));
    SLE \b6_OKctIF[155]  (.D(b4_nUAi[308]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[309]));
    SLE \b6_OKctIF[416]  (.D(b4_nUAi[47]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[48]));
    SLE \b6_OKctIF[97]  (.D(b4_nUAi[366]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[367]));
    SLE \b6_OKctIF[272]  (.D(b4_nUAi[191]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[192]));
    SLE \b6_OKctIF[142]  (.D(b4_nUAi[321]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[322]));
    SLE \b6_OKctIF[79]  (.D(b4_nUAi[384]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[385]));
    SLE \b6_OKctIF[294]  (.D(b4_nUAi[169]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[170]));
    SLE \b6_OKctIF[10]  (.D(b4_nUAi[453]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[454]));
    SLE \b6_OKctIF[96]  (.D(b4_nUAi[367]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[368]));
    SLE \b6_OKctIF[93]  (.D(b4_nUAi[370]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[371]));
    SLE \b6_OKctIF[62]  (.D(b4_nUAi[401]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[402]));
    SLE \b6_OKctIF[237]  (.D(b4_nUAi[226]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[227]));
    SLE \b6_OKctIF[119]  (.D(b4_nUAi[344]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[345]));
    SLE \b6_OKctIF[219]  (.D(b4_nUAi[244]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[245]));
    SLE \b6_OKctIF[69]  (.D(b4_nUAi[394]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[395]));
    SLE \b6_OKctIF[305]  (.D(b4_nUAi[158]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[159]));
    SLE \b6_OKctIF[205]  (.D(b4_nUAi[258]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[259]));
    SLE \b6_OKctIF[385]  (.D(b4_nUAi[78]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[79]));
    SLE \b6_OKctIF[307]  (.D(b4_nUAi[156]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[157]));
    SLE \b6_OKctIF[285]  (.D(b4_nUAi[178]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[179]));
    SLE \b6_OKctIF[387]  (.D(b4_nUAi[76]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[77]));
    SLE \b6_OKctIF[372]  (.D(b4_nUAi[91]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[92]));
    SLE \b6_OKctIF[298]  (.D(b4_nUAi[165]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[166]));
    SLE \b6_OKctIF[224]  (.D(b4_nUAi[239]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[240]));
    SLE \b6_OKctIF[210]  (.D(b4_nUAi[253]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[254]));
    SLE \b6_OKctIF[115]  (.D(b4_nUAi[348]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[349]));
    SLE \b6_OKctIF[0]  (.D(b4_nUAi[463]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b7_PSyi3wy));
    SLE \b6_OKctIF[84]  (.D(b4_nUAi[379]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[380]));
    SLE \b6_OKctIF[176]  (.D(b4_nUAi[287]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[288]));
    SLE \b6_OKctIF[70]  (.D(b4_nUAi[393]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[394]));
    SLE \b6_OKctIF[364]  (.D(b4_nUAi[99]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[100]));
    SLE \b6_OKctIF[228]  (.D(b4_nUAi[235]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[236]));
    SLE \b6_OKctIF[60]  (.D(b4_nUAi[403]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[404]));
    SLE \b6_OKctIF[425]  (.D(b4_nUAi[38]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[39]));
    SLE \b6_OKctIF[81]  (.D(b4_nUAi[382]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[383]));
    SLE \b6_OKctIF[462]  (.D(b4_nUAi[1]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[2]));
    SLE \b6_OKctIF[271]  (.D(b4_nUAi[192]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[193]));
    SLE \b6_OKctIF[232]  (.D(b4_nUAi[231]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[232]));
    SLE \b6_OKctIF[92]  (.D(b4_nUAi[371]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[372]));
    SLE \b6_OKctIF[444]  (.D(b4_nUAi[19]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[20]));
    SLE \b6_OKctIF[99]  (.D(b4_nUAi[364]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[365]));
    SLE \b6_OKctIF[87]  (.D(b4_nUAi[376]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[377]));
    SLE \b6_OKctIF[429]  (.D(b4_nUAi[34]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[35]));
    SLE \b6_OKctIF[190]  (.D(b4_nUAi[273]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[274]));
    SLE \b6_OKctIF[86]  (.D(b4_nUAi[377]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[378]));
    SLE \b6_OKctIF[83]  (.D(b4_nUAi[380]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[381]));
    SLE \b6_OKctIF[332]  (.D(b4_nUAi[131]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[132]));
    SLE \b6_OKctIF[254]  (.D(b4_nUAi[209]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[210]));
    SLE \b6_OKctIF[421]  (.D(b4_nUAi[42]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[43]));
    SLE \b6_OKctIF[193]  (.D(b4_nUAi[270]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[271]));
    SLE \b6_OKctIF[136]  (.D(b4_nUAi[327]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[328]));
    SLE \b6_OKctIF[120]  (.D(b4_nUAi[343]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[344]));
    SLE \b6_OKctIF[423]  (.D(b4_nUAi[40]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[41]));
    SLE \b6_OKctIF[258]  (.D(b4_nUAi[205]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[206]));
    SLE \b6_OKctIF[90]  (.D(b4_nUAi[373]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[374]));
    SLE \b6_OKctIF[247]  (.D(b4_nUAi[216]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[217]));
    SLE \b6_OKctIF[455]  (.D(b4_nUAi[8]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[9]));
    SLE \b6_OKctIF[192]  (.D(b4_nUAi[271]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[272]));
    SLE \b6_OKctIF[123]  (.D(b4_nUAi[340]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[341]));
    SLE \b6_OKctIF[108]  (.D(b4_nUAi[355]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[356]));
    SLE \b6_OKctIF[365]  (.D(b4_nUAi[98]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[99]));
    SLE \b6_OKctIF[265]  (.D(b4_nUAi[198]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[199]));
    SLE \b6_OKctIF[188]  (.D(b4_nUAi[275]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[276]));
    SLE \b6_OKctIF[367]  (.D(b4_nUAi[96]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[97]));
    SLE \b6_OKctIF[48]  (.D(b4_nUAi[415]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[416]));
    SLE \b6_OKctIF[45]  (.D(b4_nUAi[418]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[419]));
    SLE \b6_OKctIF[231]  (.D(b4_nUAi[232]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[233]));
    SLE \b6_OKctIF[214]  (.D(b4_nUAi[249]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[250]));
    SLE \b6_OKctIF[459]  (.D(b4_nUAi[4]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[5]));
    SLE \b6_OKctIF[122]  (.D(b4_nUAi[341]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[342]));
    SLE \b6_OKctIF[82]  (.D(b4_nUAi[381]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[382]));
    SLE \b6_OKctIF[218]  (.D(b4_nUAi[245]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[246]));
    SLE \b6_OKctIF[89]  (.D(b4_nUAi[374]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[375]));
    SLE \b6_OKctIF[415]  (.D(b4_nUAi[48]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[49]));
    SLE \b6_OKctIF[451]  (.D(b4_nUAi[12]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[13]));
    SLE \b6_OKctIF[203]  (.D(b4_nUAi[260]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[261]));
    SLE \b6_OKctIF[150]  (.D(b4_nUAi[313]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[314]));
    SLE \b6_OKctIF[283]  (.D(b4_nUAi[180]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[181]));
    SLE \b6_OKctIF[242]  (.D(b4_nUAi[221]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[222]));
    SLE \b6_OKctIF[453]  (.D(b4_nUAi[10]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[11]));
    SLE \b6_OKctIF[303]  (.D(b4_nUAi[160]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[161]));
    SLE \b6_OKctIF[383]  (.D(b4_nUAi[80]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[81]));
    SLE \b6_OKctIF[419]  (.D(b4_nUAi[44]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[45]));
    SLE \b6_OKctIF[306]  (.D(b4_nUAi[157]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[158]));
    SLE \b6_OKctIF[153]  (.D(b4_nUAi[310]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[311]));
    SLE \b6_OKctIF[101]  (.D(b4_nUAi[362]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[363]));
    SLE \b6_OKctIF[386]  (.D(b4_nUAi[77]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[78]));
    SLE \b6_OKctIF[181]  (.D(b4_nUAi[282]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[283]));
    SLE \b6_OKctIF[80]  (.D(b4_nUAi[383]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[384]));
    SLE \b6_OKctIF[1]  (.D(b4_nUAi[462]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[463]));
    SLE \b6_OKctIF[342]  (.D(b4_nUAi[121]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[122]));
    SLE \b6_OKctIF[174]  (.D(b4_nUAi[289]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[290]));
    SLE \b6_OKctIF[411]  (.D(b4_nUAi[52]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[53]));
    SLE \b6_OKctIF[152]  (.D(b4_nUAi[311]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[312]));
    SLE \b6_OKctIF[146]  (.D(b4_nUAi[317]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[318]));
    SLE \b6_OKctIF[110]  (.D(b4_nUAi[353]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[354]));
    SLE \b6_OKctIF[370]  (.D(b4_nUAi[93]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[94]));
    SLE \b6_OKctIF[413]  (.D(b4_nUAi[50]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[51]));
    SLE \b6_OKctIF[424]  (.D(b4_nUAi[39]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[40]));
    SLE \b6_OKctIF[177]  (.D(b4_nUAi[286]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[287]));
    SLE \b6_OKctIF[113]  (.D(b4_nUAi[350]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[351]));
    SLE \b6_OKctIF[438]  (.D(b4_nUAi[25]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[26]));
    SLE \b6_OKctIF[168]  (.D(b4_nUAi[295]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[296]));
    SLE \b6_OKctIF[297]  (.D(b4_nUAi[166]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[167]));
    SLE \b6_OKctIF[241]  (.D(b4_nUAi[222]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[223]));
    SLE \b6_OKctIF[112]  (.D(b4_nUAi[351]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[352]));
    SLE \b6_OKctIF[227]  (.D(b4_nUAi[236]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[237]));
    SLE \b6_OKctIF[276]  (.D(b4_nUAi[187]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[188]));
    SLE \b6_OKctIF[134]  (.D(b4_nUAi[329]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[330]));
    SLE \b6_OKctIF[309]  (.D(b4_nUAi[154]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[155]));
    SLE \b6_OKctIF[389]  (.D(b4_nUAi[74]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[75]));
    SLE \b6_OKctIF[406]  (.D(b4_nUAi[57]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[58]));
    SLE \b6_OKctIF[330]  (.D(b4_nUAi[133]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[134]));
    SLE \b6_OKctIF[263]  (.D(b4_nUAi[200]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[201]));
    SLE \b6_OKctIF[454]  (.D(b4_nUAi[9]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[10]));
    SLE \b6_OKctIF[363]  (.D(b4_nUAi[100]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[101]));
    SLE \b6_OKctIF[109]  (.D(b4_nUAi[354]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[355]));
    SLE \b6_OKctIF[209]  (.D(b4_nUAi[254]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[255]));
    SLE \b6_OKctIF[189]  (.D(b4_nUAi[274]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[275]));
    SLE \b6_OKctIF[292]  (.D(b4_nUAi[171]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[172]));
    SLE \b6_OKctIF[289]  (.D(b4_nUAi[174]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[175]));
    SLE \b6_OKctIF[137]  (.D(b4_nUAi[326]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[327]));
    SLE \b6_OKctIF[366]  (.D(b4_nUAi[97]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[98]));
    SLE \b6_OKctIF[161]  (.D(b4_nUAi[302]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[303]));
    SLE \b6_OKctIF[8]  (.D(b4_nUAi[455]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[456]));
    SLE \b6_OKctIF[200]  (.D(b4_nUAi[263]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[264]));
    SLE \b6_OKctIF[371]  (.D(b4_nUAi[92]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[93]));
    SLE \b6_OKctIF[280]  (.D(b4_nUAi[183]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[184]));
    SLE \b6_OKctIF[105]  (.D(b4_nUAi[358]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[359]));
    SLE \b6_OKctIF[185]  (.D(b4_nUAi[278]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[279]));
    SLE \b6_OKctIF[392]  (.D(b4_nUAi[71]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[72]));
    SLE \b6_OKctIF[378]  (.D(b4_nUAi[85]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[86]));
    SLE \b6_OKctIF[222]  (.D(b4_nUAi[241]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[242]));
    SLE \b6_OKctIF[414]  (.D(b4_nUAi[49]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[50]));
    SLE \b6_OKctIF[257]  (.D(b4_nUAi[206]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[207]));
    SLE \b6_OKctIF[236]  (.D(b4_nUAi[227]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[228]));
    SLE \b6_OKctIF[196]  (.D(b4_nUAi[267]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[268]));
    SLE \b6_OKctIF[448]  (.D(b4_nUAi[15]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[16]));
    SLE \b6_OKctIF[322]  (.D(b4_nUAi[141]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[142]));
    SLE \b6_OKctIF[28]  (.D(b4_nUAi[435]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[436]));
    SLE \b6_OKctIF[25]  (.D(b4_nUAi[438]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[439]));
    SLE \b6_OKctIF[126]  (.D(b4_nUAi[337]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[338]));
    SLE \b6_OKctIF[291]  (.D(b4_nUAi[172]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[173]));
    SLE \b6_OKctIF[217]  (.D(b4_nUAi[246]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[247]));
    SLE \b6_OKctIF[144]  (.D(b4_nUAi[319]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[320]));
    SLE \b6_OKctIF[44]  (.D(b4_nUAi[419]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[420]));
    SLE \b6_OKctIF[369]  (.D(b4_nUAi[94]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[95]));
    SLE \b6_OKctIF[331]  (.D(b4_nUAi[132]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[133]));
    SLE \b6_OKctIF[252]  (.D(b4_nUAi[211]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[212]));
    SLE \b6_OKctIF[340]  (.D(b4_nUAi[123]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[124]));
    SLE \b6_OKctIF[338]  (.D(b4_nUAi[125]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[126]));
    SLE \b6_OKctIF[221]  (.D(b4_nUAi[242]), .CLK(IICE_comm2iice[11]), 
        .EN(b6_OKctIF4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_nUAi[243]));
    
endmodule


module b8_1LbcQDr1_x_26_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [128:128] mdiclink_reg;
input  [26:26] b11_OFWNT9L_8tZ;
input  [385:384] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[128]), .B(
        b11_OFWNT9L_8tZ[26]), .C(b4_nUAi[385]), .D(b4_nUAi[384]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[128]), .B(
        b11_OFWNT9L_8tZ[26]), .C(b4_nUAi[385]), .D(b4_nUAi[384]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_80_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [74:74] mdiclink_reg;
input  [80:80] b11_OFWNT9L_8tZ;
input  [223:222] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[74]), .B(
        b11_OFWNT9L_8tZ[80]), .C(b4_nUAi[223]), .D(b4_nUAi[222]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[74]), .B(
        b11_OFWNT9L_8tZ[80]), .C(b4_nUAi[223]), .D(b4_nUAi[222]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_3_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [151:151] mdiclink_reg;
input  [3:3] b11_OFWNT9L_8tZ;
input  [454:453] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[151]), .B(
        b11_OFWNT9L_8tZ[3]), .C(b4_nUAi[454]), .D(b4_nUAi[453]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[151]), .B(
        b11_OFWNT9L_8tZ[3]), .C(b4_nUAi[454]), .D(b4_nUAi[453]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_27_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [127:127] mdiclink_reg;
input  [27:27] b11_OFWNT9L_8tZ;
input  [383:381] b4_nUAi;
output [127:127] b6_2ZTGIf;

    wire b3_P_F_6_bm_39, b3_P_F_6_am_39, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_39), .B(
        b4_nUAi[383]), .C(b3_P_F_6_am_39), .Y(b6_2ZTGIf[127]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[127]), .B(
        b11_OFWNT9L_8tZ[27]), .C(b4_nUAi[382]), .D(b4_nUAi[381]), .Y(
        b3_P_F_6_am_39));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[127]), .B(
        b11_OFWNT9L_8tZ[27]), .C(b4_nUAi[381]), .D(b4_nUAi[382]), .Y(
        b3_P_F_6_bm_39));
    
endmodule


module b8_1LbcQDr1_x_140_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [14:14] mdiclink_reg;
input  [140:140] b11_OFWNT9L_8tZ;
input  [44:42] b4_nUAi;
output [14:14] b6_2ZTGIf;

    wire b3_P_F_6_bm_67, b3_P_F_6_am_67, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_67), .B(
        b4_nUAi[44]), .C(b3_P_F_6_am_67), .Y(b6_2ZTGIf[14]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[14]), .B(
        b11_OFWNT9L_8tZ[140]), .C(b4_nUAi[43]), .D(b4_nUAi[42]), .Y(
        b3_P_F_6_am_67));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[14]), .B(
        b11_OFWNT9L_8tZ[140]), .C(b4_nUAi[42]), .D(b4_nUAi[43]), .Y(
        b3_P_F_6_bm_67));
    
endmodule


module b8_1LbcQDr1_x_83_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [71:71] mdiclink_reg;
input  [83:83] b11_OFWNT9L_8tZ;
input  [215:213] b4_nUAi;
output [71:71] b6_2ZTGIf;

    wire b3_P_F_6_bm_15, b3_P_F_6_am_15, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_15), .B(
        b4_nUAi[215]), .C(b3_P_F_6_am_15), .Y(b6_2ZTGIf[71]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[71]), .B(
        b11_OFWNT9L_8tZ[83]), .C(b4_nUAi[214]), .D(b4_nUAi[213]), .Y(
        b3_P_F_6_am_15));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[71]), .B(
        b11_OFWNT9L_8tZ[83]), .C(b4_nUAi[213]), .D(b4_nUAi[214]), .Y(
        b3_P_F_6_bm_15));
    
endmodule


module b8_1LbcQDr1_x_143_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [11:11] mdiclink_reg;
input  [143:143] b11_OFWNT9L_8tZ;
input  [35:33] b4_nUAi;
output [11:11] b6_2ZTGIf;

    wire b3_P_F_6_bm_70, b3_P_F_6_am_70, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_70), .B(
        b4_nUAi[35]), .C(b3_P_F_6_am_70), .Y(b6_2ZTGIf[11]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[11]), .B(
        b11_OFWNT9L_8tZ[143]), .C(b4_nUAi[34]), .D(b4_nUAi[33]), .Y(
        b3_P_F_6_am_70));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[11]), .B(
        b11_OFWNT9L_8tZ[143]), .C(b4_nUAi[33]), .D(b4_nUAi[34]), .Y(
        b3_P_F_6_bm_70));
    
endmodule


module b8_1LbcQDr1_x_34_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [120:120] mdiclink_reg;
input  [34:34] b11_OFWNT9L_8tZ;
input  [361:360] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[120]), .B(
        b11_OFWNT9L_8tZ[34]), .C(b4_nUAi[361]), .D(b4_nUAi[360]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[120]), .B(
        b11_OFWNT9L_8tZ[34]), .C(b4_nUAi[361]), .D(b4_nUAi[360]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_84_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [70:70] mdiclink_reg;
input  [84:84] b11_OFWNT9L_8tZ;
input  [212:210] b4_nUAi;
output [70:70] b6_2ZTGIf;

    wire b3_P_F_6_bm_16, b3_P_F_6_am_16, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_16), .B(
        b4_nUAi[212]), .C(b3_P_F_6_am_16), .Y(b6_2ZTGIf[70]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[70]), .B(
        b11_OFWNT9L_8tZ[84]), .C(b4_nUAi[211]), .D(b4_nUAi[210]), .Y(
        b3_P_F_6_am_16));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[70]), .B(
        b11_OFWNT9L_8tZ[84]), .C(b4_nUAi[210]), .D(b4_nUAi[211]), .Y(
        b3_P_F_6_bm_16));
    
endmodule


module b8_1LbcQDr1_x_144_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [10:10] mdiclink_reg;
input  [144:144] b11_OFWNT9L_8tZ;
input  [31:30] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[10]), .B(
        b11_OFWNT9L_8tZ[144]), .C(b4_nUAi[31]), .D(b4_nUAi[30]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[10]), .B(
        b11_OFWNT9L_8tZ[144]), .C(b4_nUAi[31]), .D(b4_nUAi[30]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_103_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [51:51] mdiclink_reg;
input  [103:103] b11_OFWNT9L_8tZ;
input  [154:153] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[51]), .B(
        b11_OFWNT9L_8tZ[103]), .C(b4_nUAi[154]), .D(b4_nUAi[153]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[51]), .B(
        b11_OFWNT9L_8tZ[103]), .C(b4_nUAi[154]), .D(b4_nUAi[153]), .Y(
        N_25));
    
endmodule


module b9_O2yyf_fG2_x_8_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [5:5] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[5]));
    
endmodule


module b9_O2yyf_fG2_x_5_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [8:8] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[8]));
    
endmodule


module b9_O2yyf_fG2_x_4_0(
       b13_CZS0wfY_d_FH9,
       b6_2ZTGIf_1,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_10,
       b6_2ZTGIf_9,
       b6_2ZTGIf_8,
       b6_2ZTGIf_0,
       b4_nUAi_0,
       b4_nUAi_6,
       b4_nUAi_12,
       b4_nUAi_15,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2
    );
output [9:9] b13_CZS0wfY_d_FH9;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_0;
input  b4_nUAi_0;
input  b4_nUAi_6;
input  b4_nUAi_12;
input  b4_nUAi_15;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;

    wire o_2_net_1, o_1_net_1, o_0_net_1, o_7_net_1, o_5_net_1, 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_1), .D(N_27), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_0), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_3), .D(N_27_0), .Y(o_1_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8000) )  o_7 (.A(b6_2ZTGIf_10), .B(b6_2ZTGIf_9), 
        .C(b6_2ZTGIf_8), .D(b6_2ZTGIf_0), .Y(o_7_net_1));
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_1), .B(b4_nUAi_12), .C(
        b6_2ZTGIf_5), .D(N_27_1), .Y(o_0_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_2_net_1), .B(o_1_net_1), .C(
        o_7_net_1), .D(o_5_net_1), .Y(b13_CZS0wfY_d_FH9[9]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25_2), .B(b4_nUAi_15), .C(
        o_0_net_1), .D(N_27_2), .Y(o_5_net_1));
    
endmodule


module b9_O2yyf_fG2_x_13_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [0:0] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[0]));
    
endmodule


module b9_O2yyf_fG2_x_9_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [4:4] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[4]));
    
endmodule


module b9_O2yyf_fG2_x_10_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [3:3] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[3]));
    
endmodule


module b9_O2yyf_fG2_x_11_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [2:2] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[2]));
    
endmodule


module b9_O2yyf_fG2_x_6_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [7:7] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[7]));
    
endmodule


module b9_O2yyf_fG2_x_0_0(
       b14_CZS0wfY_d_FH9m,
       b11_uUT0JC4gFrY
    );
input  [9:0] b14_CZS0wfY_d_FH9m;
output [1:1] b11_uUT0JC4gFrY;

    wire o_6_net_1, o_5_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h8000) )  o_6 (.A(b14_CZS0wfY_d_FH9m[3]), .B(
        b14_CZS0wfY_d_FH9m[2]), .C(b14_CZS0wfY_d_FH9m[1]), .D(
        b14_CZS0wfY_d_FH9m[0]), .Y(o_6_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(b14_CZS0wfY_d_FH9m[9]), .B(
        b14_CZS0wfY_d_FH9m[8]), .C(o_6_net_1), .D(o_5_net_1), .Y(
        b11_uUT0JC4gFrY[1]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h8000) )  o_5 (.A(b14_CZS0wfY_d_FH9m[7]), .B(
        b14_CZS0wfY_d_FH9m[6]), .C(b14_CZS0wfY_d_FH9m[5]), .D(
        b14_CZS0wfY_d_FH9m[4]), .Y(o_5_net_1));
    
endmodule


module b9_O2yyf_fG2_x_12_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [1:1] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[1]));
    
endmodule


module b9_O2yyf_fG2_x_7_0(
       b13_CZS0wfY_d_FH9,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4
    );
output [6:6] b13_CZS0wfY_d_FH9;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;

    wire o_5_net_1, o_4_net_1, o_3_net_1, o_2_net_1, o_1_net_1, 
        o_0_net_1, o_11_net_1, o_12_net_1, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hE020) )  o_0 (.A(N_25_4), .B(b4_nUAi_9), .C(
        b6_2ZTGIf_10), .D(N_27_4), .Y(o_0_net_1));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hE020) )  o_3 (.A(N_25_1), .B(b4_nUAi_0), .C(
        b6_2ZTGIf_7), .D(N_27_1), .Y(o_3_net_1));
    CFG4 #( .INIT(16'h8000) )  o_11 (.A(b6_2ZTGIf_11), .B(b6_2ZTGIf_2), 
        .C(b6_2ZTGIf_1), .D(b6_2ZTGIf_0), .Y(o_11_net_1));
    CFG4 #( .INIT(16'hE020) )  o_1 (.A(N_25_3), .B(b4_nUAi_6), .C(
        b6_2ZTGIf_9), .D(N_27_3), .Y(o_1_net_1));
    CFG4 #( .INIT(16'hE020) )  o_2 (.A(N_25_2), .B(b4_nUAi_3), .C(
        b6_2ZTGIf_8), .D(N_27_2), .Y(o_2_net_1));
    CFG4 #( .INIT(16'hE020) )  o_5 (.A(N_25), .B(b4_nUAi_24), .C(
        b6_2ZTGIf_3), .D(N_27), .Y(o_5_net_1));
    CFG4 #( .INIT(16'hE020) )  o_4 (.A(N_25_0), .B(b4_nUAi_30), .C(
        b6_2ZTGIf_5), .D(N_27_0), .Y(o_4_net_1));
    CFG4 #( .INIT(16'h8000) )  o_12 (.A(o_3_net_1), .B(o_2_net_1), .C(
        o_1_net_1), .D(o_0_net_1), .Y(o_12_net_1));
    CFG4 #( .INIT(16'h8000) )  o (.A(o_4_net_1), .B(o_5_net_1), .C(
        o_12_net_1), .D(o_11_net_1), .Y(b13_CZS0wfY_d_FH9[6]));
    
endmodule


module b16_CRGcTCua_eH4_uui_x_0(
       b11_uUT0JC4gFrY,
       b6_2ZTGIf_3,
       b6_2ZTGIf_5,
       b6_2ZTGIf_7,
       b6_2ZTGIf_8,
       b6_2ZTGIf_9,
       b6_2ZTGIf_10,
       b6_2ZTGIf_11,
       b6_2ZTGIf_2,
       b6_2ZTGIf_1,
       b6_2ZTGIf_0,
       b6_2ZTGIf_19,
       b6_2ZTGIf_21,
       b6_2ZTGIf_23,
       b6_2ZTGIf_24,
       b6_2ZTGIf_25,
       b6_2ZTGIf_26,
       b6_2ZTGIf_27,
       b6_2ZTGIf_18,
       b6_2ZTGIf_17,
       b6_2ZTGIf_16,
       b6_2ZTGIf_35,
       b6_2ZTGIf_37,
       b6_2ZTGIf_39,
       b6_2ZTGIf_40,
       b6_2ZTGIf_41,
       b6_2ZTGIf_42,
       b6_2ZTGIf_43,
       b6_2ZTGIf_34,
       b6_2ZTGIf_33,
       b6_2ZTGIf_32,
       b6_2ZTGIf_51,
       b6_2ZTGIf_53,
       b6_2ZTGIf_55,
       b6_2ZTGIf_56,
       b6_2ZTGIf_57,
       b6_2ZTGIf_58,
       b6_2ZTGIf_59,
       b6_2ZTGIf_50,
       b6_2ZTGIf_49,
       b6_2ZTGIf_48,
       b6_2ZTGIf_67,
       b6_2ZTGIf_69,
       b6_2ZTGIf_71,
       b6_2ZTGIf_72,
       b6_2ZTGIf_73,
       b6_2ZTGIf_74,
       b6_2ZTGIf_75,
       b6_2ZTGIf_66,
       b6_2ZTGIf_65,
       b6_2ZTGIf_64,
       b6_2ZTGIf_83,
       b6_2ZTGIf_85,
       b6_2ZTGIf_87,
       b6_2ZTGIf_88,
       b6_2ZTGIf_89,
       b6_2ZTGIf_90,
       b6_2ZTGIf_91,
       b6_2ZTGIf_82,
       b6_2ZTGIf_81,
       b6_2ZTGIf_80,
       b6_2ZTGIf_99,
       b6_2ZTGIf_101,
       b6_2ZTGIf_103,
       b6_2ZTGIf_104,
       b6_2ZTGIf_105,
       b6_2ZTGIf_106,
       b6_2ZTGIf_107,
       b6_2ZTGIf_98,
       b6_2ZTGIf_97,
       b6_2ZTGIf_96,
       b6_2ZTGIf_115,
       b6_2ZTGIf_117,
       b6_2ZTGIf_119,
       b6_2ZTGIf_120,
       b6_2ZTGIf_121,
       b6_2ZTGIf_122,
       b6_2ZTGIf_123,
       b6_2ZTGIf_114,
       b6_2ZTGIf_113,
       b6_2ZTGIf_112,
       b6_2ZTGIf_131,
       b6_2ZTGIf_133,
       b6_2ZTGIf_135,
       b6_2ZTGIf_136,
       b6_2ZTGIf_137,
       b6_2ZTGIf_138,
       b6_2ZTGIf_139,
       b6_2ZTGIf_130,
       b6_2ZTGIf_129,
       b6_2ZTGIf_128,
       b6_2ZTGIf_141,
       b6_2ZTGIf_143,
       b6_2ZTGIf_145,
       b6_2ZTGIf_150,
       b6_2ZTGIf_149,
       b6_2ZTGIf_148,
       b6_2ZTGIf_140,
       b4_nUAi_24,
       b4_nUAi_30,
       b4_nUAi_0,
       b4_nUAi_3,
       b4_nUAi_6,
       b4_nUAi_9,
       b4_nUAi_72,
       b4_nUAi_78,
       b4_nUAi_48,
       b4_nUAi_51,
       b4_nUAi_54,
       b4_nUAi_57,
       b4_nUAi_120,
       b4_nUAi_126,
       b4_nUAi_96,
       b4_nUAi_99,
       b4_nUAi_102,
       b4_nUAi_105,
       b4_nUAi_168,
       b4_nUAi_174,
       b4_nUAi_144,
       b4_nUAi_147,
       b4_nUAi_150,
       b4_nUAi_153,
       b4_nUAi_216,
       b4_nUAi_222,
       b4_nUAi_192,
       b4_nUAi_195,
       b4_nUAi_198,
       b4_nUAi_201,
       b4_nUAi_264,
       b4_nUAi_270,
       b4_nUAi_240,
       b4_nUAi_243,
       b4_nUAi_246,
       b4_nUAi_249,
       b4_nUAi_312,
       b4_nUAi_318,
       b4_nUAi_288,
       b4_nUAi_291,
       b4_nUAi_294,
       b4_nUAi_297,
       b4_nUAi_360,
       b4_nUAi_366,
       b4_nUAi_336,
       b4_nUAi_339,
       b4_nUAi_342,
       b4_nUAi_345,
       b4_nUAi_408,
       b4_nUAi_414,
       b4_nUAi_384,
       b4_nUAi_387,
       b4_nUAi_390,
       b4_nUAi_393,
       b4_nUAi_438,
       b4_nUAi_444,
       b4_nUAi_450,
       b4_nUAi_453,
       BW_clk_c,
       N_25,
       N_27,
       N_25_0,
       N_27_0,
       N_25_1,
       N_27_1,
       N_25_2,
       N_27_2,
       N_25_3,
       N_27_3,
       N_25_4,
       N_27_4,
       N_25_5,
       N_27_5,
       N_25_6,
       N_27_6,
       N_25_7,
       N_27_7,
       N_25_8,
       N_27_8,
       N_25_9,
       N_27_9,
       N_25_10,
       N_27_10,
       N_25_11,
       N_27_11,
       N_25_12,
       N_27_12,
       N_25_13,
       N_27_13,
       N_25_14,
       N_27_14,
       N_25_15,
       N_27_15,
       N_25_16,
       N_27_16,
       N_25_17,
       N_27_17,
       N_25_18,
       N_27_18,
       N_25_19,
       N_27_19,
       N_25_20,
       N_27_20,
       N_25_21,
       N_27_21,
       N_25_22,
       N_27_22,
       N_25_23,
       N_27_23,
       N_25_24,
       N_27_24,
       N_25_25,
       N_27_25,
       N_25_26,
       N_27_26,
       N_25_27,
       N_27_27,
       N_25_28,
       N_27_28,
       N_25_29,
       N_27_29,
       N_25_30,
       N_27_30,
       N_25_31,
       N_27_31,
       N_25_32,
       N_27_32,
       N_25_33,
       N_27_33,
       N_25_34,
       N_27_34,
       N_25_35,
       N_27_35,
       N_25_36,
       N_27_36,
       N_25_37,
       N_27_37,
       N_25_38,
       N_27_38,
       N_25_39,
       N_27_39,
       N_25_40,
       N_27_40,
       N_25_41,
       N_27_41,
       N_25_42,
       N_27_42,
       N_25_43,
       N_27_43,
       N_25_44,
       N_27_44,
       N_25_45,
       N_27_45,
       N_25_46,
       N_27_46,
       N_25_47,
       N_27_47,
       N_25_48,
       N_27_48,
       N_25_49,
       N_27_49,
       N_25_50,
       N_27_50,
       N_25_51,
       N_27_51,
       N_25_52,
       N_27_52,
       N_25_53,
       N_27_53,
       N_25_54,
       N_27_54,
       N_25_55,
       N_27_55,
       N_25_56,
       N_27_56
    );
output [1:1] b11_uUT0JC4gFrY;
input  b6_2ZTGIf_3;
input  b6_2ZTGIf_5;
input  b6_2ZTGIf_7;
input  b6_2ZTGIf_8;
input  b6_2ZTGIf_9;
input  b6_2ZTGIf_10;
input  b6_2ZTGIf_11;
input  b6_2ZTGIf_2;
input  b6_2ZTGIf_1;
input  b6_2ZTGIf_0;
input  b6_2ZTGIf_19;
input  b6_2ZTGIf_21;
input  b6_2ZTGIf_23;
input  b6_2ZTGIf_24;
input  b6_2ZTGIf_25;
input  b6_2ZTGIf_26;
input  b6_2ZTGIf_27;
input  b6_2ZTGIf_18;
input  b6_2ZTGIf_17;
input  b6_2ZTGIf_16;
input  b6_2ZTGIf_35;
input  b6_2ZTGIf_37;
input  b6_2ZTGIf_39;
input  b6_2ZTGIf_40;
input  b6_2ZTGIf_41;
input  b6_2ZTGIf_42;
input  b6_2ZTGIf_43;
input  b6_2ZTGIf_34;
input  b6_2ZTGIf_33;
input  b6_2ZTGIf_32;
input  b6_2ZTGIf_51;
input  b6_2ZTGIf_53;
input  b6_2ZTGIf_55;
input  b6_2ZTGIf_56;
input  b6_2ZTGIf_57;
input  b6_2ZTGIf_58;
input  b6_2ZTGIf_59;
input  b6_2ZTGIf_50;
input  b6_2ZTGIf_49;
input  b6_2ZTGIf_48;
input  b6_2ZTGIf_67;
input  b6_2ZTGIf_69;
input  b6_2ZTGIf_71;
input  b6_2ZTGIf_72;
input  b6_2ZTGIf_73;
input  b6_2ZTGIf_74;
input  b6_2ZTGIf_75;
input  b6_2ZTGIf_66;
input  b6_2ZTGIf_65;
input  b6_2ZTGIf_64;
input  b6_2ZTGIf_83;
input  b6_2ZTGIf_85;
input  b6_2ZTGIf_87;
input  b6_2ZTGIf_88;
input  b6_2ZTGIf_89;
input  b6_2ZTGIf_90;
input  b6_2ZTGIf_91;
input  b6_2ZTGIf_82;
input  b6_2ZTGIf_81;
input  b6_2ZTGIf_80;
input  b6_2ZTGIf_99;
input  b6_2ZTGIf_101;
input  b6_2ZTGIf_103;
input  b6_2ZTGIf_104;
input  b6_2ZTGIf_105;
input  b6_2ZTGIf_106;
input  b6_2ZTGIf_107;
input  b6_2ZTGIf_98;
input  b6_2ZTGIf_97;
input  b6_2ZTGIf_96;
input  b6_2ZTGIf_115;
input  b6_2ZTGIf_117;
input  b6_2ZTGIf_119;
input  b6_2ZTGIf_120;
input  b6_2ZTGIf_121;
input  b6_2ZTGIf_122;
input  b6_2ZTGIf_123;
input  b6_2ZTGIf_114;
input  b6_2ZTGIf_113;
input  b6_2ZTGIf_112;
input  b6_2ZTGIf_131;
input  b6_2ZTGIf_133;
input  b6_2ZTGIf_135;
input  b6_2ZTGIf_136;
input  b6_2ZTGIf_137;
input  b6_2ZTGIf_138;
input  b6_2ZTGIf_139;
input  b6_2ZTGIf_130;
input  b6_2ZTGIf_129;
input  b6_2ZTGIf_128;
input  b6_2ZTGIf_141;
input  b6_2ZTGIf_143;
input  b6_2ZTGIf_145;
input  b6_2ZTGIf_150;
input  b6_2ZTGIf_149;
input  b6_2ZTGIf_148;
input  b6_2ZTGIf_140;
input  b4_nUAi_24;
input  b4_nUAi_30;
input  b4_nUAi_0;
input  b4_nUAi_3;
input  b4_nUAi_6;
input  b4_nUAi_9;
input  b4_nUAi_72;
input  b4_nUAi_78;
input  b4_nUAi_48;
input  b4_nUAi_51;
input  b4_nUAi_54;
input  b4_nUAi_57;
input  b4_nUAi_120;
input  b4_nUAi_126;
input  b4_nUAi_96;
input  b4_nUAi_99;
input  b4_nUAi_102;
input  b4_nUAi_105;
input  b4_nUAi_168;
input  b4_nUAi_174;
input  b4_nUAi_144;
input  b4_nUAi_147;
input  b4_nUAi_150;
input  b4_nUAi_153;
input  b4_nUAi_216;
input  b4_nUAi_222;
input  b4_nUAi_192;
input  b4_nUAi_195;
input  b4_nUAi_198;
input  b4_nUAi_201;
input  b4_nUAi_264;
input  b4_nUAi_270;
input  b4_nUAi_240;
input  b4_nUAi_243;
input  b4_nUAi_246;
input  b4_nUAi_249;
input  b4_nUAi_312;
input  b4_nUAi_318;
input  b4_nUAi_288;
input  b4_nUAi_291;
input  b4_nUAi_294;
input  b4_nUAi_297;
input  b4_nUAi_360;
input  b4_nUAi_366;
input  b4_nUAi_336;
input  b4_nUAi_339;
input  b4_nUAi_342;
input  b4_nUAi_345;
input  b4_nUAi_408;
input  b4_nUAi_414;
input  b4_nUAi_384;
input  b4_nUAi_387;
input  b4_nUAi_390;
input  b4_nUAi_393;
input  b4_nUAi_438;
input  b4_nUAi_444;
input  b4_nUAi_450;
input  b4_nUAi_453;
input  BW_clk_c;
input  N_25;
input  N_27;
input  N_25_0;
input  N_27_0;
input  N_25_1;
input  N_27_1;
input  N_25_2;
input  N_27_2;
input  N_25_3;
input  N_27_3;
input  N_25_4;
input  N_27_4;
input  N_25_5;
input  N_27_5;
input  N_25_6;
input  N_27_6;
input  N_25_7;
input  N_27_7;
input  N_25_8;
input  N_27_8;
input  N_25_9;
input  N_27_9;
input  N_25_10;
input  N_27_10;
input  N_25_11;
input  N_27_11;
input  N_25_12;
input  N_27_12;
input  N_25_13;
input  N_27_13;
input  N_25_14;
input  N_27_14;
input  N_25_15;
input  N_27_15;
input  N_25_16;
input  N_27_16;
input  N_25_17;
input  N_27_17;
input  N_25_18;
input  N_27_18;
input  N_25_19;
input  N_27_19;
input  N_25_20;
input  N_27_20;
input  N_25_21;
input  N_27_21;
input  N_25_22;
input  N_27_22;
input  N_25_23;
input  N_27_23;
input  N_25_24;
input  N_27_24;
input  N_25_25;
input  N_27_25;
input  N_25_26;
input  N_27_26;
input  N_25_27;
input  N_27_27;
input  N_25_28;
input  N_27_28;
input  N_25_29;
input  N_27_29;
input  N_25_30;
input  N_27_30;
input  N_25_31;
input  N_27_31;
input  N_25_32;
input  N_27_32;
input  N_25_33;
input  N_27_33;
input  N_25_34;
input  N_27_34;
input  N_25_35;
input  N_27_35;
input  N_25_36;
input  N_27_36;
input  N_25_37;
input  N_27_37;
input  N_25_38;
input  N_27_38;
input  N_25_39;
input  N_27_39;
input  N_25_40;
input  N_27_40;
input  N_25_41;
input  N_27_41;
input  N_25_42;
input  N_27_42;
input  N_25_43;
input  N_27_43;
input  N_25_44;
input  N_27_44;
input  N_25_45;
input  N_27_45;
input  N_25_46;
input  N_27_46;
input  N_25_47;
input  N_27_47;
input  N_25_48;
input  N_27_48;
input  N_25_49;
input  N_27_49;
input  N_25_50;
input  N_27_50;
input  N_25_51;
input  N_27_51;
input  N_25_52;
input  N_27_52;
input  N_25_53;
input  N_27_53;
input  N_25_54;
input  N_27_54;
input  N_25_55;
input  N_27_55;
input  N_25_56;
input  N_27_56;

    wire \b14_CZS0wfY_d_FH9m[9]_net_1 , VCC_net_1, 
        \b13_CZS0wfY_d_FH9[9] , GND_net_1, 
        \b14_CZS0wfY_d_FH9m[8]_net_1 , \b13_CZS0wfY_d_FH9[8] , 
        \b14_CZS0wfY_d_FH9m[7]_net_1 , \b13_CZS0wfY_d_FH9[7] , 
        \b14_CZS0wfY_d_FH9m[6]_net_1 , \b13_CZS0wfY_d_FH9[6] , 
        \b14_CZS0wfY_d_FH9m[5]_net_1 , \b13_CZS0wfY_d_FH9[5] , 
        \b14_CZS0wfY_d_FH9m[4]_net_1 , \b13_CZS0wfY_d_FH9[4] , 
        \b14_CZS0wfY_d_FH9m[3]_net_1 , \b13_CZS0wfY_d_FH9[3] , 
        \b14_CZS0wfY_d_FH9m[2]_net_1 , \b13_CZS0wfY_d_FH9[2] , 
        \b14_CZS0wfY_d_FH9m[1]_net_1 , \b13_CZS0wfY_d_FH9[1] , 
        \b14_CZS0wfY_d_FH9m[0]_net_1 , \b13_CZS0wfY_d_FH9[0] ;
    
    b9_O2yyf_fG2_x_8_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_c (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[5] }), .b4_nUAi_24(
        b4_nUAi_264), .b4_nUAi_30(b4_nUAi_270), .b4_nUAi_0(b4_nUAi_240)
        , .b4_nUAi_3(b4_nUAi_243), .b4_nUAi_6(b4_nUAi_246), .b4_nUAi_9(
        b4_nUAi_249), .b6_2ZTGIf_3(b6_2ZTGIf_83), .b6_2ZTGIf_5(
        b6_2ZTGIf_85), .b6_2ZTGIf_7(b6_2ZTGIf_87), .b6_2ZTGIf_8(
        b6_2ZTGIf_88), .b6_2ZTGIf_9(b6_2ZTGIf_89), .b6_2ZTGIf_10(
        b6_2ZTGIf_90), .b6_2ZTGIf_11(b6_2ZTGIf_91), .b6_2ZTGIf_2(
        b6_2ZTGIf_82), .b6_2ZTGIf_1(b6_2ZTGIf_81), .b6_2ZTGIf_0(
        b6_2ZTGIf_80), .N_25(N_25_29), .N_27(N_27_29), .N_25_0(N_25_30)
        , .N_27_0(N_27_30), .N_25_1(N_25_31), .N_27_1(N_27_31), 
        .N_25_2(N_25_32), .N_27_2(N_27_32), .N_25_3(N_25_33), .N_27_3(
        N_27_33), .N_25_4(N_25_34), .N_27_4(N_27_34));
    b9_O2yyf_fG2_x_5_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_F (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[8] }), .b4_nUAi_24(
        b4_nUAi_408), .b4_nUAi_30(b4_nUAi_414), .b4_nUAi_0(b4_nUAi_384)
        , .b4_nUAi_3(b4_nUAi_387), .b4_nUAi_6(b4_nUAi_390), .b4_nUAi_9(
        b4_nUAi_393), .b6_2ZTGIf_3(b6_2ZTGIf_131), .b6_2ZTGIf_5(
        b6_2ZTGIf_133), .b6_2ZTGIf_7(b6_2ZTGIf_135), .b6_2ZTGIf_8(
        b6_2ZTGIf_136), .b6_2ZTGIf_9(b6_2ZTGIf_137), .b6_2ZTGIf_10(
        b6_2ZTGIf_138), .b6_2ZTGIf_11(b6_2ZTGIf_139), .b6_2ZTGIf_2(
        b6_2ZTGIf_130), .b6_2ZTGIf_1(b6_2ZTGIf_129), .b6_2ZTGIf_0(
        b6_2ZTGIf_128), .N_25(N_25_47), .N_27(N_27_47), .N_25_0(
        N_25_48), .N_27_0(N_27_48), .N_25_1(N_25_49), .N_27_1(N_27_49), 
        .N_25_2(N_25_50), .N_27_2(N_27_50), .N_25_3(N_25_51), .N_27_3(
        N_27_51), .N_25_4(N_25_52), .N_27_4(N_27_52));
    b9_O2yyf_fG2_x_4_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_d (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[9] }), .b6_2ZTGIf_1(
        b6_2ZTGIf_141), .b6_2ZTGIf_3(b6_2ZTGIf_143), .b6_2ZTGIf_5(
        b6_2ZTGIf_145), .b6_2ZTGIf_10(b6_2ZTGIf_150), .b6_2ZTGIf_9(
        b6_2ZTGIf_149), .b6_2ZTGIf_8(b6_2ZTGIf_148), .b6_2ZTGIf_0(
        b6_2ZTGIf_140), .b4_nUAi_0(b4_nUAi_438), .b4_nUAi_6(
        b4_nUAi_444), .b4_nUAi_12(b4_nUAi_450), .b4_nUAi_15(
        b4_nUAi_453), .N_25(N_25_53), .N_27(N_27_53), .N_25_0(N_25_54), 
        .N_27_0(N_27_54), .N_25_1(N_25_55), .N_27_1(N_27_55), .N_25_2(
        N_25_56), .N_27_2(N_27_56));
    SLE \b14_CZS0wfY_d_FH9m[4]  (.D(\b13_CZS0wfY_d_FH9[4] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[4]_net_1 ));
    b9_O2yyf_fG2_x_13_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_9 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[0] }), .b4_nUAi_24(
        b4_nUAi_24), .b4_nUAi_30(b4_nUAi_30), .b4_nUAi_0(b4_nUAi_0), 
        .b4_nUAi_3(b4_nUAi_3), .b4_nUAi_6(b4_nUAi_6), .b4_nUAi_9(
        b4_nUAi_9), .b6_2ZTGIf_3(b6_2ZTGIf_3), .b6_2ZTGIf_5(
        b6_2ZTGIf_5), .b6_2ZTGIf_7(b6_2ZTGIf_7), .b6_2ZTGIf_8(
        b6_2ZTGIf_8), .b6_2ZTGIf_9(b6_2ZTGIf_9), .b6_2ZTGIf_10(
        b6_2ZTGIf_10), .b6_2ZTGIf_11(b6_2ZTGIf_11), .b6_2ZTGIf_2(
        b6_2ZTGIf_2), .b6_2ZTGIf_1(b6_2ZTGIf_1), .b6_2ZTGIf_0(
        b6_2ZTGIf_0), .N_25(N_25), .N_27(N_27), .N_25_0(N_25_0), 
        .N_27_0(N_27_0), .N_25_1(N_25_1), .N_27_1(N_27_1), .N_25_2(
        N_25_2), .N_27_2(N_27_2), .N_25_3(N_25_3), .N_27_3(N_27_3), 
        .N_25_4(N_25_4), .N_27_4(N_27_4));
    GND GND (.Y(GND_net_1));
    b9_O2yyf_fG2_x_9_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_8 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[4] }), .b4_nUAi_24(
        b4_nUAi_216), .b4_nUAi_30(b4_nUAi_222), .b4_nUAi_0(b4_nUAi_192)
        , .b4_nUAi_3(b4_nUAi_195), .b4_nUAi_6(b4_nUAi_198), .b4_nUAi_9(
        b4_nUAi_201), .b6_2ZTGIf_3(b6_2ZTGIf_67), .b6_2ZTGIf_5(
        b6_2ZTGIf_69), .b6_2ZTGIf_7(b6_2ZTGIf_71), .b6_2ZTGIf_8(
        b6_2ZTGIf_72), .b6_2ZTGIf_9(b6_2ZTGIf_73), .b6_2ZTGIf_10(
        b6_2ZTGIf_74), .b6_2ZTGIf_11(b6_2ZTGIf_75), .b6_2ZTGIf_2(
        b6_2ZTGIf_66), .b6_2ZTGIf_1(b6_2ZTGIf_65), .b6_2ZTGIf_0(
        b6_2ZTGIf_64), .N_25(N_25_23), .N_27(N_27_23), .N_25_0(N_25_24)
        , .N_27_0(N_27_24), .N_25_1(N_25_25), .N_27_1(N_27_25), 
        .N_25_2(N_25_26), .N_27_2(N_27_26), .N_25_3(N_25_27), .N_27_3(
        N_27_27), .N_25_4(N_25_28), .N_27_4(N_27_28));
    b9_O2yyf_fG2_x_10_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_I (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[3] }), .b4_nUAi_24(
        b4_nUAi_168), .b4_nUAi_30(b4_nUAi_174), .b4_nUAi_0(b4_nUAi_144)
        , .b4_nUAi_3(b4_nUAi_147), .b4_nUAi_6(b4_nUAi_150), .b4_nUAi_9(
        b4_nUAi_153), .b6_2ZTGIf_3(b6_2ZTGIf_51), .b6_2ZTGIf_5(
        b6_2ZTGIf_53), .b6_2ZTGIf_7(b6_2ZTGIf_55), .b6_2ZTGIf_8(
        b6_2ZTGIf_56), .b6_2ZTGIf_9(b6_2ZTGIf_57), .b6_2ZTGIf_10(
        b6_2ZTGIf_58), .b6_2ZTGIf_11(b6_2ZTGIf_59), .b6_2ZTGIf_2(
        b6_2ZTGIf_50), .b6_2ZTGIf_1(b6_2ZTGIf_49), .b6_2ZTGIf_0(
        b6_2ZTGIf_48), .N_25(N_25_17), .N_27(N_27_17), .N_25_0(N_25_18)
        , .N_27_0(N_27_18), .N_25_1(N_25_19), .N_27_1(N_27_19), 
        .N_25_2(N_25_20), .N_27_2(N_27_20), .N_25_3(N_25_21), .N_27_3(
        N_27_21), .N_25_4(N_25_22), .N_27_4(N_27_22));
    SLE \b14_CZS0wfY_d_FH9m[3]  (.D(\b13_CZS0wfY_d_FH9[3] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[3]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[1]  (.D(\b13_CZS0wfY_d_FH9[1] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[1]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[5]  (.D(\b13_CZS0wfY_d_FH9[5] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[5]_net_1 ));
    b9_O2yyf_fG2_x_11_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_0 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[2] }), .b4_nUAi_24(
        b4_nUAi_120), .b4_nUAi_30(b4_nUAi_126), .b4_nUAi_0(b4_nUAi_96), 
        .b4_nUAi_3(b4_nUAi_99), .b4_nUAi_6(b4_nUAi_102), .b4_nUAi_9(
        b4_nUAi_105), .b6_2ZTGIf_3(b6_2ZTGIf_35), .b6_2ZTGIf_5(
        b6_2ZTGIf_37), .b6_2ZTGIf_7(b6_2ZTGIf_39), .b6_2ZTGIf_8(
        b6_2ZTGIf_40), .b6_2ZTGIf_9(b6_2ZTGIf_41), .b6_2ZTGIf_10(
        b6_2ZTGIf_42), .b6_2ZTGIf_11(b6_2ZTGIf_43), .b6_2ZTGIf_2(
        b6_2ZTGIf_34), .b6_2ZTGIf_1(b6_2ZTGIf_33), .b6_2ZTGIf_0(
        b6_2ZTGIf_32), .N_25(N_25_11), .N_27(N_27_11), .N_25_0(N_25_12)
        , .N_27_0(N_27_12), .N_25_1(N_25_13), .N_27_1(N_27_13), 
        .N_25_2(N_25_14), .N_27_2(N_27_14), .N_25_3(N_25_15), .N_27_3(
        N_27_15), .N_25_4(N_25_16), .N_27_4(N_27_16));
    SLE \b14_CZS0wfY_d_FH9m[6]  (.D(\b13_CZS0wfY_d_FH9[6] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[6]_net_1 ));
    b9_O2yyf_fG2_x_6_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_1 (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[7] }), .b4_nUAi_24(
        b4_nUAi_360), .b4_nUAi_30(b4_nUAi_366), .b4_nUAi_0(b4_nUAi_336)
        , .b4_nUAi_3(b4_nUAi_339), .b4_nUAi_6(b4_nUAi_342), .b4_nUAi_9(
        b4_nUAi_345), .b6_2ZTGIf_3(b6_2ZTGIf_115), .b6_2ZTGIf_5(
        b6_2ZTGIf_117), .b6_2ZTGIf_7(b6_2ZTGIf_119), .b6_2ZTGIf_8(
        b6_2ZTGIf_120), .b6_2ZTGIf_9(b6_2ZTGIf_121), .b6_2ZTGIf_10(
        b6_2ZTGIf_122), .b6_2ZTGIf_11(b6_2ZTGIf_123), .b6_2ZTGIf_2(
        b6_2ZTGIf_114), .b6_2ZTGIf_1(b6_2ZTGIf_113), .b6_2ZTGIf_0(
        b6_2ZTGIf_112), .N_25(N_25_41), .N_27(N_27_41), .N_25_0(
        N_25_42), .N_27_0(N_27_42), .N_25_1(N_25_43), .N_27_1(N_27_43), 
        .N_25_2(N_25_44), .N_27_2(N_27_44), .N_25_3(N_25_45), .N_27_3(
        N_27_45), .N_25_4(N_25_46), .N_27_4(N_27_46));
    SLE \b14_CZS0wfY_d_FH9m[9]  (.D(\b13_CZS0wfY_d_FH9[9] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[9]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[7]  (.D(\b13_CZS0wfY_d_FH9[7] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[7]_net_1 ));
    b9_O2yyf_fG2_x_0_0 b25_O2yyf_fG2_MiQA1E6_Z_lnxob (
        .b14_CZS0wfY_d_FH9m({\b14_CZS0wfY_d_FH9m[9]_net_1 , 
        \b14_CZS0wfY_d_FH9m[8]_net_1 , \b14_CZS0wfY_d_FH9m[7]_net_1 , 
        \b14_CZS0wfY_d_FH9m[6]_net_1 , \b14_CZS0wfY_d_FH9m[5]_net_1 , 
        \b14_CZS0wfY_d_FH9m[4]_net_1 , \b14_CZS0wfY_d_FH9m[3]_net_1 , 
        \b14_CZS0wfY_d_FH9m[2]_net_1 , \b14_CZS0wfY_d_FH9m[1]_net_1 , 
        \b14_CZS0wfY_d_FH9m[0]_net_1 }), .b11_uUT0JC4gFrY({
        b11_uUT0JC4gFrY[1]}));
    SLE \b14_CZS0wfY_d_FH9m[2]  (.D(\b13_CZS0wfY_d_FH9[2] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[2]_net_1 ));
    SLE \b14_CZS0wfY_d_FH9m[0]  (.D(\b13_CZS0wfY_d_FH9[0] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    b9_O2yyf_fG2_x_12_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_a (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[1] }), .b4_nUAi_24(
        b4_nUAi_72), .b4_nUAi_30(b4_nUAi_78), .b4_nUAi_0(b4_nUAi_48), 
        .b4_nUAi_3(b4_nUAi_51), .b4_nUAi_6(b4_nUAi_54), .b4_nUAi_9(
        b4_nUAi_57), .b6_2ZTGIf_3(b6_2ZTGIf_19), .b6_2ZTGIf_5(
        b6_2ZTGIf_21), .b6_2ZTGIf_7(b6_2ZTGIf_23), .b6_2ZTGIf_8(
        b6_2ZTGIf_24), .b6_2ZTGIf_9(b6_2ZTGIf_25), .b6_2ZTGIf_10(
        b6_2ZTGIf_26), .b6_2ZTGIf_11(b6_2ZTGIf_27), .b6_2ZTGIf_2(
        b6_2ZTGIf_18), .b6_2ZTGIf_1(b6_2ZTGIf_17), .b6_2ZTGIf_0(
        b6_2ZTGIf_16), .N_25(N_25_5), .N_27(N_27_5), .N_25_0(N_25_6), 
        .N_27_0(N_27_6), .N_25_1(N_25_7), .N_27_1(N_27_7), .N_25_2(
        N_25_8), .N_27_2(N_27_8), .N_25_3(N_25_9), .N_27_3(N_27_9), 
        .N_25_4(N_25_10), .N_27_4(N_27_10));
    b9_O2yyf_fG2_x_7_0 b27_O2yyf_fG2_MiQA1E6_r_lnxob_S (
        .b13_CZS0wfY_d_FH9({\b13_CZS0wfY_d_FH9[6] }), .b4_nUAi_24(
        b4_nUAi_312), .b4_nUAi_30(b4_nUAi_318), .b4_nUAi_0(b4_nUAi_288)
        , .b4_nUAi_3(b4_nUAi_291), .b4_nUAi_6(b4_nUAi_294), .b4_nUAi_9(
        b4_nUAi_297), .b6_2ZTGIf_3(b6_2ZTGIf_99), .b6_2ZTGIf_5(
        b6_2ZTGIf_101), .b6_2ZTGIf_7(b6_2ZTGIf_103), .b6_2ZTGIf_8(
        b6_2ZTGIf_104), .b6_2ZTGIf_9(b6_2ZTGIf_105), .b6_2ZTGIf_10(
        b6_2ZTGIf_106), .b6_2ZTGIf_11(b6_2ZTGIf_107), .b6_2ZTGIf_2(
        b6_2ZTGIf_98), .b6_2ZTGIf_1(b6_2ZTGIf_97), .b6_2ZTGIf_0(
        b6_2ZTGIf_96), .N_25(N_25_35), .N_27(N_27_35), .N_25_0(N_25_36)
        , .N_27_0(N_27_36), .N_25_1(N_25_37), .N_27_1(N_27_37), 
        .N_25_2(N_25_38), .N_27_2(N_27_38), .N_25_3(N_25_39), .N_27_3(
        N_27_39), .N_25_4(N_25_40), .N_27_4(N_27_40));
    SLE \b14_CZS0wfY_d_FH9m[8]  (.D(\b13_CZS0wfY_d_FH9[8] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b14_CZS0wfY_d_FH9m[8]_net_1 ));
    
endmodule


module b8_1LbcQDr1_x_104_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [50:50] mdiclink_reg;
input  [104:104] b11_OFWNT9L_8tZ;
input  [151:150] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[50]), .B(
        b11_OFWNT9L_8tZ[104]), .C(b4_nUAi[151]), .D(b4_nUAi[150]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[50]), .B(
        b11_OFWNT9L_8tZ[104]), .C(b4_nUAi[151]), .D(b4_nUAi[150]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_72_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [82:82] mdiclink_reg;
input  [72:72] b11_OFWNT9L_8tZ;
input  [247:246] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[82]), .B(
        b11_OFWNT9L_8tZ[72]), .C(b4_nUAi[247]), .D(b4_nUAi[246]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[82]), .B(
        b11_OFWNT9L_8tZ[72]), .C(b4_nUAi[247]), .D(b4_nUAi[246]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_33_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [121:121] mdiclink_reg;
input  [33:33] b11_OFWNT9L_8tZ;
input  [365:363] b4_nUAi;
output [121:121] b6_2ZTGIf;

    wire b3_P_F_6_bm_44, b3_P_F_6_am_44, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_44), .B(
        b4_nUAi[365]), .C(b3_P_F_6_am_44), .Y(b6_2ZTGIf[121]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[121]), .B(
        b11_OFWNT9L_8tZ[33]), .C(b4_nUAi[364]), .D(b4_nUAi[363]), .Y(
        b3_P_F_6_am_44));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[121]), .B(
        b11_OFWNT9L_8tZ[33]), .C(b4_nUAi[363]), .D(b4_nUAi[364]), .Y(
        b3_P_F_6_bm_44));
    
endmodule


module b8_1LbcQDr1_x_129_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [25:25] mdiclink_reg;
input  [129:129] b11_OFWNT9L_8tZ;
input  [77:75] b4_nUAi;
output [25:25] b6_2ZTGIf;

    wire b3_P_F_6_bm_81, b3_P_F_6_am_81, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_81), .B(
        b4_nUAi[77]), .C(b3_P_F_6_am_81), .Y(b6_2ZTGIf[25]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[25]), .B(
        b11_OFWNT9L_8tZ[129]), .C(b4_nUAi[76]), .D(b4_nUAi[75]), .Y(
        b3_P_F_6_am_81));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[25]), .B(
        b11_OFWNT9L_8tZ[129]), .C(b4_nUAi[75]), .D(b4_nUAi[76]), .Y(
        b3_P_F_6_bm_81));
    
endmodule


module b8_1LbcQDr1_x_89_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [65:65] mdiclink_reg;
input  [89:89] b11_OFWNT9L_8tZ;
input  [196:195] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[65]), .B(
        b11_OFWNT9L_8tZ[89]), .C(b4_nUAi[196]), .D(b4_nUAi[195]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[65]), .B(
        b11_OFWNT9L_8tZ[89]), .C(b4_nUAi[196]), .D(b4_nUAi[195]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_120_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [34:34] mdiclink_reg;
input  [120:120] b11_OFWNT9L_8tZ;
input  [103:102] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[34]), .B(
        b11_OFWNT9L_8tZ[120]), .C(b4_nUAi[103]), .D(b4_nUAi[102]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[34]), .B(
        b11_OFWNT9L_8tZ[120]), .C(b4_nUAi[103]), .D(b4_nUAi[102]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_90_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [64:64] mdiclink_reg;
input  [90:90] b11_OFWNT9L_8tZ;
input  [193:192] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[64]), .B(
        b11_OFWNT9L_8tZ[90]), .C(b4_nUAi[193]), .D(b4_nUAi[192]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[64]), .B(
        b11_OFWNT9L_8tZ[90]), .C(b4_nUAi[193]), .D(b4_nUAi[192]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_10_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [144:144] mdiclink_reg;
input  [10:10] b11_OFWNT9L_8tZ;
input  [434:432] b4_nUAi;
output [144:144] b6_2ZTGIf;

    wire b3_P_F_6_bm_65, b3_P_F_6_am_65, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_65), .B(
        b4_nUAi[434]), .C(b3_P_F_6_am_65), .Y(b6_2ZTGIf[144]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[144]), .B(
        b11_OFWNT9L_8tZ[10]), .C(b4_nUAi[433]), .D(b4_nUAi[432]), .Y(
        b3_P_F_6_am_65));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[144]), .B(
        b11_OFWNT9L_8tZ[10]), .C(b4_nUAi[432]), .D(b4_nUAi[433]), .Y(
        b3_P_F_6_bm_65));
    
endmodule


module b8_1LbcQDr1_x_8_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [146:146] mdiclink_reg;
input  [8:8] b11_OFWNT9L_8tZ;
input  [439:438] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[146]), .B(
        b11_OFWNT9L_8tZ[8]), .C(b4_nUAi[439]), .D(b4_nUAi[438]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[146]), .B(
        b11_OFWNT9L_8tZ[8]), .C(b4_nUAi[439]), .D(b4_nUAi[438]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_1_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [153:153] mdiclink_reg;
input  [1:1] b11_OFWNT9L_8tZ;
input  [461:459] b4_nUAi;
output [153:153] b6_2ZTGIf;

    wire b3_P_F_6_bm_60, b3_P_F_6_am_60, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_60), .B(
        b4_nUAi[461]), .C(b3_P_F_6_am_60), .Y(b6_2ZTGIf[153]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[153]), .B(
        b11_OFWNT9L_8tZ[1]), .C(b4_nUAi[460]), .D(b4_nUAi[459]), .Y(
        b3_P_F_6_am_60));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[153]), .B(
        b11_OFWNT9L_8tZ[1]), .C(b4_nUAi[459]), .D(b4_nUAi[460]), .Y(
        b3_P_F_6_bm_60));
    
endmodule


module b8_1LbcQDr1_x_130_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [24:24] mdiclink_reg;
input  [130:130] b11_OFWNT9L_8tZ;
input  [73:72] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[24]), .B(
        b11_OFWNT9L_8tZ[130]), .C(b4_nUAi[73]), .D(b4_nUAi[72]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[24]), .B(
        b11_OFWNT9L_8tZ[130]), .C(b4_nUAi[73]), .D(b4_nUAi[72]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_132_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [22:22] mdiclink_reg;
input  [132:132] b11_OFWNT9L_8tZ;
input  [68:66] b4_nUAi;
output [22:22] b6_2ZTGIf;

    wire b3_P_F_6_bm_83, b3_P_F_6_am_83, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_83), .B(
        b4_nUAi[68]), .C(b3_P_F_6_am_83), .Y(b6_2ZTGIf[22]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[22]), .B(
        b11_OFWNT9L_8tZ[132]), .C(b4_nUAi[67]), .D(b4_nUAi[66]), .Y(
        b3_P_F_6_am_83));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[22]), .B(
        b11_OFWNT9L_8tZ[132]), .C(b4_nUAi[66]), .D(b4_nUAi[67]), .Y(
        b3_P_F_6_bm_83));
    
endmodule


module b8_1LbcQDr1_x_92_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [62:62] mdiclink_reg;
input  [92:92] b11_OFWNT9L_8tZ;
input  [188:186] b4_nUAi;
output [62:62] b6_2ZTGIf;

    wire b3_P_F_6_bm_0, b3_P_F_6_am_0, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_0), .B(
        b4_nUAi[188]), .C(b3_P_F_6_am_0), .Y(b6_2ZTGIf[62]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[62]), .B(
        b11_OFWNT9L_8tZ[92]), .C(b4_nUAi[187]), .D(b4_nUAi[186]), .Y(
        b3_P_F_6_am_0));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[62]), .B(
        b11_OFWNT9L_8tZ[92]), .C(b4_nUAi[186]), .D(b4_nUAi[187]), .Y(
        b3_P_F_6_bm_0));
    
endmodule


module b8_1LbcQDr1_x_113_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [41:41] mdiclink_reg;
input  [113:113] b11_OFWNT9L_8tZ;
input  [125:123] b4_nUAi;
output [41:41] b6_2ZTGIf;

    wire b3_P_F_6_bm_91, b3_P_F_6_am_91, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_91), .B(
        b4_nUAi[125]), .C(b3_P_F_6_am_91), .Y(b6_2ZTGIf[41]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[41]), .B(
        b11_OFWNT9L_8tZ[113]), .C(b4_nUAi[124]), .D(b4_nUAi[123]), .Y(
        b3_P_F_6_am_91));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[41]), .B(
        b11_OFWNT9L_8tZ[113]), .C(b4_nUAi[123]), .D(b4_nUAi[124]), .Y(
        b3_P_F_6_bm_91));
    
endmodule


module b8_1LbcQDr1_x_76_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [78:78] mdiclink_reg;
input  [76:76] b11_OFWNT9L_8tZ;
input  [236:234] b4_nUAi;
output [78:78] b6_2ZTGIf;

    wire b3_P_F_6_bm_10, b3_P_F_6_am_10, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_10), .B(
        b4_nUAi[236]), .C(b3_P_F_6_am_10), .Y(b6_2ZTGIf[78]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[78]), .B(
        b11_OFWNT9L_8tZ[76]), .C(b4_nUAi[235]), .D(b4_nUAi[234]), .Y(
        b3_P_F_6_am_10));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[78]), .B(
        b11_OFWNT9L_8tZ[76]), .C(b4_nUAi[234]), .D(b4_nUAi[235]), .Y(
        b3_P_F_6_bm_10));
    
endmodule


module b8_1LbcQDr1_x_136_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [18:18] mdiclink_reg;
input  [136:136] b11_OFWNT9L_8tZ;
input  [55:54] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[18]), .B(
        b11_OFWNT9L_8tZ[136]), .C(b4_nUAi[55]), .D(b4_nUAi[54]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[18]), .B(
        b11_OFWNT9L_8tZ[136]), .C(b4_nUAi[55]), .D(b4_nUAi[54]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_67_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [87:87] mdiclink_reg;
input  [67:67] b11_OFWNT9L_8tZ;
input  [263:261] b4_nUAi;
output [87:87] b6_2ZTGIf;

    wire b3_P_F_6_bm_25, b3_P_F_6_am_25, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_25), .B(
        b4_nUAi[263]), .C(b3_P_F_6_am_25), .Y(b6_2ZTGIf[87]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[87]), .B(
        b11_OFWNT9L_8tZ[67]), .C(b4_nUAi[262]), .D(b4_nUAi[261]), .Y(
        b3_P_F_6_am_25));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[87]), .B(
        b11_OFWNT9L_8tZ[67]), .C(b4_nUAi[261]), .D(b4_nUAi[262]), .Y(
        b3_P_F_6_bm_25));
    
endmodule


module b8_1LbcQDr1_x_114_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [40:40] mdiclink_reg;
input  [114:114] b11_OFWNT9L_8tZ;
input  [121:120] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[40]), .B(
        b11_OFWNT9L_8tZ[114]), .C(b4_nUAi[121]), .D(b4_nUAi[120]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[40]), .B(
        b11_OFWNT9L_8tZ[114]), .C(b4_nUAi[121]), .D(b4_nUAi[120]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_118_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [36:36] mdiclink_reg;
input  [118:118] b11_OFWNT9L_8tZ;
input  [110:108] b4_nUAi;
output [36:36] b6_2ZTGIf;

    wire b3_P_F_6_bm_95, b3_P_F_6_am_95, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_95), .B(
        b4_nUAi[110]), .C(b3_P_F_6_am_95), .Y(b6_2ZTGIf[36]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[36]), .B(
        b11_OFWNT9L_8tZ[118]), .C(b4_nUAi[109]), .D(b4_nUAi[108]), .Y(
        b3_P_F_6_am_95));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[36]), .B(
        b11_OFWNT9L_8tZ[118]), .C(b4_nUAi[108]), .D(b4_nUAi[109]), .Y(
        b3_P_F_6_bm_95));
    
endmodule


module b8_1LbcQDr1_x_96_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [58:58] mdiclink_reg;
input  [96:96] b11_OFWNT9L_8tZ;
input  [175:174] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[58]), .B(
        b11_OFWNT9L_8tZ[96]), .C(b4_nUAi[175]), .D(b4_nUAi[174]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[58]), .B(
        b11_OFWNT9L_8tZ[96]), .C(b4_nUAi[175]), .D(b4_nUAi[174]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_31_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [123:123] mdiclink_reg;
input  [31:31] b11_OFWNT9L_8tZ;
input  [371:369] b4_nUAi;
output [123:123] b6_2ZTGIf;

    wire b3_P_F_6_bm_43, b3_P_F_6_am_43, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_43), .B(
        b4_nUAi[371]), .C(b3_P_F_6_am_43), .Y(b6_2ZTGIf[123]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[123]), .B(
        b11_OFWNT9L_8tZ[31]), .C(b4_nUAi[370]), .D(b4_nUAi[369]), .Y(
        b3_P_F_6_am_43));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[123]), .B(
        b11_OFWNT9L_8tZ[31]), .C(b4_nUAi[369]), .D(b4_nUAi[370]), .Y(
        b3_P_F_6_bm_43));
    
endmodule


module b8_1LbcQDr1_x_75_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [79:79] mdiclink_reg;
input  [75:75] b11_OFWNT9L_8tZ;
input  [239:237] b4_nUAi;
output [79:79] b6_2ZTGIf;

    wire b3_P_F_6_bm_9, b3_P_F_6_am_9, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_9), .B(
        b4_nUAi[239]), .C(b3_P_F_6_am_9), .Y(b6_2ZTGIf[79]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[79]), .B(
        b11_OFWNT9L_8tZ[75]), .C(b4_nUAi[238]), .D(b4_nUAi[237]), .Y(
        b3_P_F_6_am_9));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[79]), .B(
        b11_OFWNT9L_8tZ[75]), .C(b4_nUAi[237]), .D(b4_nUAi[238]), .Y(
        b3_P_F_6_bm_9));
    
endmodule


module b8_1LbcQDr1_x_135_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [19:19] mdiclink_reg;
input  [135:135] b11_OFWNT9L_8tZ;
input  [58:57] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[19]), .B(
        b11_OFWNT9L_8tZ[135]), .C(b4_nUAi[58]), .D(b4_nUAi[57]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[19]), .B(
        b11_OFWNT9L_8tZ[135]), .C(b4_nUAi[58]), .D(b4_nUAi[57]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_20_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [134:134] mdiclink_reg;
input  [20:20] b11_OFWNT9L_8tZ;
input  [404:402] b4_nUAi;
output [134:134] b6_2ZTGIf;

    wire b3_P_F_6_bm_56, b3_P_F_6_am_56, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_56), .B(
        b4_nUAi[404]), .C(b3_P_F_6_am_56), .Y(b6_2ZTGIf[134]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[134]), .B(
        b11_OFWNT9L_8tZ[20]), .C(b4_nUAi[403]), .D(b4_nUAi[402]), .Y(
        b3_P_F_6_am_56));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[134]), .B(
        b11_OFWNT9L_8tZ[20]), .C(b4_nUAi[402]), .D(b4_nUAi[403]), .Y(
        b3_P_F_6_bm_56));
    
endmodule


module b8_1LbcQDr1_x_95_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [59:59] mdiclink_reg;
input  [95:95] b11_OFWNT9L_8tZ;
input  [179:177] b4_nUAi;
output [59:59] b6_2ZTGIf;

    wire b3_P_F_6_bm_3, b3_P_F_6_am_3, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_3), .B(
        b4_nUAi[179]), .C(b3_P_F_6_am_3), .Y(b6_2ZTGIf[59]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[59]), .B(
        b11_OFWNT9L_8tZ[95]), .C(b4_nUAi[178]), .D(b4_nUAi[177]), .Y(
        b3_P_F_6_am_3));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[59]), .B(
        b11_OFWNT9L_8tZ[95]), .C(b4_nUAi[177]), .D(b4_nUAi[178]), .Y(
        b3_P_F_6_bm_3));
    
endmodule


module b8_1LbcQDr1_x_150_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [4:4] mdiclink_reg;
input  [150:150] b11_OFWNT9L_8tZ;
input  [14:12] b4_nUAi;
output [4:4] b6_2ZTGIf;

    wire b3_P_F_6_bm_75, b3_P_F_6_am_75, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_75), .B(
        b4_nUAi[14]), .C(b3_P_F_6_am_75), .Y(b6_2ZTGIf[4]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[4]), .B(
        b11_OFWNT9L_8tZ[150]), .C(b4_nUAi[13]), .D(b4_nUAi[12]), .Y(
        b3_P_F_6_am_75));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[4]), .B(
        b11_OFWNT9L_8tZ[150]), .C(b4_nUAi[12]), .D(b4_nUAi[13]), .Y(
        b3_P_F_6_bm_75));
    
endmodule


module b8_1LbcQDr1_x_18_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [136:136] mdiclink_reg;
input  [18:18] b11_OFWNT9L_8tZ;
input  [409:408] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[136]), .B(
        b11_OFWNT9L_8tZ[18]), .C(b4_nUAi[409]), .D(b4_nUAi[408]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[136]), .B(
        b11_OFWNT9L_8tZ[18]), .C(b4_nUAi[409]), .D(b4_nUAi[408]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_127_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [27:27] mdiclink_reg;
input  [127:127] b11_OFWNT9L_8tZ;
input  [83:81] b4_nUAi;
output [27:27] b6_2ZTGIf;

    wire b3_P_F_6_bm_80, b3_P_F_6_am_80, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_80), .B(
        b4_nUAi[83]), .C(b3_P_F_6_am_80), .Y(b6_2ZTGIf[27]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[27]), .B(
        b11_OFWNT9L_8tZ[127]), .C(b4_nUAi[82]), .D(b4_nUAi[81]), .Y(
        b3_P_F_6_am_80));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[27]), .B(
        b11_OFWNT9L_8tZ[127]), .C(b4_nUAi[81]), .D(b4_nUAi[82]), .Y(
        b3_P_F_6_bm_80));
    
endmodule


module b8_1LbcQDr1_x_87_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [67:67] mdiclink_reg;
input  [87:87] b11_OFWNT9L_8tZ;
input  [202:201] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[67]), .B(
        b11_OFWNT9L_8tZ[87]), .C(b4_nUAi[202]), .D(b4_nUAi[201]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[67]), .B(
        b11_OFWNT9L_8tZ[87]), .C(b4_nUAi[202]), .D(b4_nUAi[201]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_40_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [114:114] mdiclink_reg;
input  [40:40] b11_OFWNT9L_8tZ;
input  [343:342] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[114]), .B(
        b11_OFWNT9L_8tZ[40]), .C(b4_nUAi[343]), .D(b4_nUAi[342]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[114]), .B(
        b11_OFWNT9L_8tZ[40]), .C(b4_nUAi[343]), .D(b4_nUAi[342]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_58_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [96:96] mdiclink_reg;
input  [58:58] b11_OFWNT9L_8tZ;
input  [289:288] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[96]), .B(
        b11_OFWNT9L_8tZ[58]), .C(b4_nUAi[289]), .D(b4_nUAi[288]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[96]), .B(
        b11_OFWNT9L_8tZ[58]), .C(b4_nUAi[289]), .D(b4_nUAi[288]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_38_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [116:116] mdiclink_reg;
input  [38:38] b11_OFWNT9L_8tZ;
input  [350:348] b4_nUAi;
output [116:116] b6_2ZTGIf;

    wire b3_P_F_6_bm_48, b3_P_F_6_am_48, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_48), .B(
        b4_nUAi[350]), .C(b3_P_F_6_am_48), .Y(b6_2ZTGIf[116]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[116]), .B(
        b11_OFWNT9L_8tZ[38]), .C(b4_nUAi[349]), .D(b4_nUAi[348]), .Y(
        b3_P_F_6_am_48));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[116]), .B(
        b11_OFWNT9L_8tZ[38]), .C(b4_nUAi[348]), .D(b4_nUAi[349]), .Y(
        b3_P_F_6_bm_48));
    
endmodule


module b8_1LbcQDr1_x_50_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [104:104] mdiclink_reg;
input  [50:50] b11_OFWNT9L_8tZ;
input  [313:312] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[104]), .B(
        b11_OFWNT9L_8tZ[50]), .C(b4_nUAi[313]), .D(b4_nUAi[312]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[104]), .B(
        b11_OFWNT9L_8tZ[50]), .C(b4_nUAi[313]), .D(b4_nUAi[312]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_121_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [33:33] mdiclink_reg;
input  [121:121] b11_OFWNT9L_8tZ;
input  [100:99] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[33]), .B(
        b11_OFWNT9L_8tZ[121]), .C(b4_nUAi[100]), .D(b4_nUAi[99]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[33]), .B(
        b11_OFWNT9L_8tZ[121]), .C(b4_nUAi[100]), .D(b4_nUAi[99]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_48_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [106:106] mdiclink_reg;
input  [48:48] b11_OFWNT9L_8tZ;
input  [319:318] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[106]), .B(
        b11_OFWNT9L_8tZ[48]), .C(b4_nUAi[319]), .D(b4_nUAi[318]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[106]), .B(
        b11_OFWNT9L_8tZ[48]), .C(b4_nUAi[319]), .D(b4_nUAi[318]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_106_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [48:48] mdiclink_reg;
input  [106:106] b11_OFWNT9L_8tZ;
input  [145:144] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[48]), .B(
        b11_OFWNT9L_8tZ[106]), .C(b4_nUAi[145]), .D(b4_nUAi[144]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[48]), .B(
        b11_OFWNT9L_8tZ[106]), .C(b4_nUAi[145]), .D(b4_nUAi[144]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_79_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [75:75] mdiclink_reg;
input  [79:79] b11_OFWNT9L_8tZ;
input  [227:225] b4_nUAi;
output [75:75] b6_2ZTGIf;

    wire b3_P_F_6_bm_13, b3_P_F_6_am_13, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_13), .B(
        b4_nUAi[227]), .C(b3_P_F_6_am_13), .Y(b6_2ZTGIf[75]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[75]), .B(
        b11_OFWNT9L_8tZ[79]), .C(b4_nUAi[226]), .D(b4_nUAi[225]), .Y(
        b3_P_F_6_am_13));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[75]), .B(
        b11_OFWNT9L_8tZ[79]), .C(b4_nUAi[225]), .D(b4_nUAi[226]), .Y(
        b3_P_F_6_bm_13));
    
endmodule


module b8_1LbcQDr1_x_139_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [15:15] mdiclink_reg;
input  [139:139] b11_OFWNT9L_8tZ;
input  [47:45] b4_nUAi;
output [15:15] b6_2ZTGIf;

    wire b3_P_F_6_bm_66, b3_P_F_6_am_66, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_66), .B(
        b4_nUAi[47]), .C(b3_P_F_6_am_66), .Y(b6_2ZTGIf[15]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[15]), .B(
        b11_OFWNT9L_8tZ[139]), .C(b4_nUAi[46]), .D(b4_nUAi[45]), .Y(
        b3_P_F_6_am_66));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[15]), .B(
        b11_OFWNT9L_8tZ[139]), .C(b4_nUAi[45]), .D(b4_nUAi[46]), .Y(
        b3_P_F_6_bm_66));
    
endmodule


module b8_1LbcQDr1_x_147_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [7:7] mdiclink_reg;
input  [147:147] b11_OFWNT9L_8tZ;
input  [23:21] b4_nUAi;
output [7:7] b6_2ZTGIf;

    wire b3_P_F_6_bm_72, b3_P_F_6_am_72, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_72), .B(
        b4_nUAi[23]), .C(b3_P_F_6_am_72), .Y(b6_2ZTGIf[7]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[7]), .B(
        b11_OFWNT9L_8tZ[147]), .C(b4_nUAi[22]), .D(b4_nUAi[21]), .Y(
        b3_P_F_6_am_72));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[7]), .B(
        b11_OFWNT9L_8tZ[147]), .C(b4_nUAi[21]), .D(b4_nUAi[22]), .Y(
        b3_P_F_6_bm_72));
    
endmodule


module b8_1LbcQDr1_x_99_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [55:55] mdiclink_reg;
input  [99:99] b11_OFWNT9L_8tZ;
input  [167:165] b4_nUAi;
output [55:55] b6_2ZTGIf;

    wire b3_P_F_6_bm_5, b3_P_F_6_am_5, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_5), .B(
        b4_nUAi[167]), .C(b3_P_F_6_am_5), .Y(b6_2ZTGIf[55]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[55]), .B(
        b11_OFWNT9L_8tZ[99]), .C(b4_nUAi[166]), .D(b4_nUAi[165]), .Y(
        b3_P_F_6_am_5));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[55]), .B(
        b11_OFWNT9L_8tZ[99]), .C(b4_nUAi[165]), .D(b4_nUAi[166]), .Y(
        b3_P_F_6_bm_5));
    
endmodule


module b8_1LbcQDr1_x_105_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [49:49] mdiclink_reg;
input  [105:105] b11_OFWNT9L_8tZ;
input  [148:147] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[49]), .B(
        b11_OFWNT9L_8tZ[105]), .C(b4_nUAi[148]), .D(b4_nUAi[147]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[49]), .B(
        b11_OFWNT9L_8tZ[105]), .C(b4_nUAi[148]), .D(b4_nUAi[147]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_110_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [44:44] mdiclink_reg;
input  [110:110] b11_OFWNT9L_8tZ;
input  [134:132] b4_nUAi;
output [44:44] b6_2ZTGIf;

    wire b3_P_F_6_bm_89, b3_P_F_6_am_89, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_89), .B(
        b4_nUAi[134]), .C(b3_P_F_6_am_89), .Y(b6_2ZTGIf[44]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[44]), .B(
        b11_OFWNT9L_8tZ[110]), .C(b4_nUAi[133]), .D(b4_nUAi[132]), .Y(
        b3_P_F_6_am_89));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[44]), .B(
        b11_OFWNT9L_8tZ[110]), .C(b4_nUAi[132]), .D(b4_nUAi[133]), .Y(
        b3_P_F_6_bm_89));
    
endmodule


module b8_1LbcQDr1_x_123_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [31:31] mdiclink_reg;
input  [123:123] b11_OFWNT9L_8tZ;
input  [95:93] b4_nUAi;
output [31:31] b6_2ZTGIf;

    wire b3_P_F_6_bm_76, b3_P_F_6_am_76, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_76), .B(
        b4_nUAi[95]), .C(b3_P_F_6_am_76), .Y(b6_2ZTGIf[31]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[31]), .B(
        b11_OFWNT9L_8tZ[123]), .C(b4_nUAi[94]), .D(b4_nUAi[93]), .Y(
        b3_P_F_6_am_76));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[31]), .B(
        b11_OFWNT9L_8tZ[123]), .C(b4_nUAi[93]), .D(b4_nUAi[94]), .Y(
        b3_P_F_6_bm_76));
    
endmodule


module b8_1LbcQDr1_x_82_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [72:72] mdiclink_reg;
input  [82:82] b11_OFWNT9L_8tZ;
input  [217:216] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[72]), .B(
        b11_OFWNT9L_8tZ[82]), .C(b4_nUAi[217]), .D(b4_nUAi[216]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[72]), .B(
        b11_OFWNT9L_8tZ[82]), .C(b4_nUAi[217]), .D(b4_nUAi[216]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_142_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [12:12] mdiclink_reg;
input  [142:142] b11_OFWNT9L_8tZ;
input  [38:36] b4_nUAi;
output [12:12] b6_2ZTGIf;

    wire b3_P_F_6_bm_69, b3_P_F_6_am_69, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_69), .B(
        b4_nUAi[38]), .C(b3_P_F_6_am_69), .Y(b6_2ZTGIf[12]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[12]), .B(
        b11_OFWNT9L_8tZ[142]), .C(b4_nUAi[37]), .D(b4_nUAi[36]), .Y(
        b3_P_F_6_am_69));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[12]), .B(
        b11_OFWNT9L_8tZ[142]), .C(b4_nUAi[36]), .D(b4_nUAi[37]), .Y(
        b3_P_F_6_bm_69));
    
endmodule


module b8_1LbcQDr1_x_124_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [30:30] mdiclink_reg;
input  [124:124] b11_OFWNT9L_8tZ;
input  [92:90] b4_nUAi;
output [30:30] b6_2ZTGIf;

    wire b3_P_F_6_bm_77, b3_P_F_6_am_77, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_77), .B(
        b4_nUAi[92]), .C(b3_P_F_6_am_77), .Y(b6_2ZTGIf[30]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[30]), .B(
        b11_OFWNT9L_8tZ[124]), .C(b4_nUAi[91]), .D(b4_nUAi[90]), .Y(
        b3_P_F_6_am_77));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[30]), .B(
        b11_OFWNT9L_8tZ[124]), .C(b4_nUAi[90]), .D(b4_nUAi[91]), .Y(
        b3_P_F_6_bm_77));
    
endmodule


module b8_1LbcQDr1_x_102_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [52:52] mdiclink_reg;
input  [102:102] b11_OFWNT9L_8tZ;
input  [158:156] b4_nUAi;
output [52:52] b6_2ZTGIf;

    wire b3_P_F_6_bm_8, b3_P_F_6_am_8, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_8), .B(
        b4_nUAi[158]), .C(b3_P_F_6_am_8), .Y(b6_2ZTGIf[52]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[52]), .B(
        b11_OFWNT9L_8tZ[102]), .C(b4_nUAi[157]), .D(b4_nUAi[156]), .Y(
        b3_P_F_6_am_8));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[52]), .B(
        b11_OFWNT9L_8tZ[102]), .C(b4_nUAi[156]), .D(b4_nUAi[157]), .Y(
        b3_P_F_6_bm_8));
    
endmodule


module b8_1LbcQDr1_x_12_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [142:142] mdiclink_reg;
input  [12:12] b11_OFWNT9L_8tZ;
input  [428:426] b4_nUAi;
output [142:142] b6_2ZTGIf;

    wire b3_P_F_6_bm_50, b3_P_F_6_am_50, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_50), .B(
        b4_nUAi[428]), .C(b3_P_F_6_am_50), .Y(b6_2ZTGIf[142]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[142]), .B(
        b11_OFWNT9L_8tZ[12]), .C(b4_nUAi[427]), .D(b4_nUAi[426]), .Y(
        b3_P_F_6_am_50));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[142]), .B(
        b11_OFWNT9L_8tZ[12]), .C(b4_nUAi[426]), .D(b4_nUAi[427]), .Y(
        b3_P_F_6_bm_50));
    
endmodule


module b8_1LbcQDr1_x_61_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [93:93] mdiclink_reg;
input  [61:61] b11_OFWNT9L_8tZ;
input  [281:279] b4_nUAi;
output [93:93] b6_2ZTGIf;

    wire b3_P_F_6_bm_21, b3_P_F_6_am_21, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_21), .B(
        b4_nUAi[281]), .C(b3_P_F_6_am_21), .Y(b6_2ZTGIf[93]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[93]), .B(
        b11_OFWNT9L_8tZ[61]), .C(b4_nUAi[280]), .D(b4_nUAi[279]), .Y(
        b3_P_F_6_am_21));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[93]), .B(
        b11_OFWNT9L_8tZ[61]), .C(b4_nUAi[279]), .D(b4_nUAi[280]), .Y(
        b3_P_F_6_bm_21));
    
endmodule


module b8_1LbcQDr1_x_148_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [6:6] mdiclink_reg;
input  [148:148] b11_OFWNT9L_8tZ;
input  [20:18] b4_nUAi;
output [6:6] b6_2ZTGIf;

    wire b3_P_F_6_bm_73, b3_P_F_6_am_73, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_73), .B(
        b4_nUAi[20]), .C(b3_P_F_6_am_73), .Y(b6_2ZTGIf[6]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[6]), .B(
        b11_OFWNT9L_8tZ[148]), .C(b4_nUAi[19]), .D(b4_nUAi[18]), .Y(
        b3_P_F_6_am_73));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[6]), .B(
        b11_OFWNT9L_8tZ[148]), .C(b4_nUAi[18]), .D(b4_nUAi[19]), .Y(
        b3_P_F_6_bm_73));
    
endmodule


module b8_1LbcQDr1_x_9_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [145:145] mdiclink_reg;
input  [9:9] b11_OFWNT9L_8tZ;
input  [437:435] b4_nUAi;
output [145:145] b6_2ZTGIf;

    wire b3_P_F_6_bm_64, b3_P_F_6_am_64, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_64), .B(
        b4_nUAi[437]), .C(b3_P_F_6_am_64), .Y(b6_2ZTGIf[145]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[145]), .B(
        b11_OFWNT9L_8tZ[9]), .C(b4_nUAi[436]), .D(b4_nUAi[435]), .Y(
        b3_P_F_6_am_64));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[145]), .B(
        b11_OFWNT9L_8tZ[9]), .C(b4_nUAi[435]), .D(b4_nUAi[436]), .Y(
        b3_P_F_6_bm_64));
    
endmodule


module b8_1LbcQDr1_x_109_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [45:45] mdiclink_reg;
input  [109:109] b11_OFWNT9L_8tZ;
input  [137:135] b4_nUAi;
output [45:45] b6_2ZTGIf;

    wire b3_P_F_6_bm_88, b3_P_F_6_am_88, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_88), .B(
        b4_nUAi[137]), .C(b3_P_F_6_am_88), .Y(b6_2ZTGIf[45]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[45]), .B(
        b11_OFWNT9L_8tZ[109]), .C(b4_nUAi[136]), .D(b4_nUAi[135]), .Y(
        b3_P_F_6_am_88));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[45]), .B(
        b11_OFWNT9L_8tZ[109]), .C(b4_nUAi[135]), .D(b4_nUAi[136]), .Y(
        b3_P_F_6_bm_88));
    
endmodule


module b8_1LbcQDr1_x_5_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [149:149] mdiclink_reg;
input  [5:5] b11_OFWNT9L_8tZ;
input  [449:447] b4_nUAi;
output [149:149] b6_2ZTGIf;

    wire b3_P_F_6_bm_62, b3_P_F_6_am_62, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_62), .B(
        b4_nUAi[449]), .C(b3_P_F_6_am_62), .Y(b6_2ZTGIf[149]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[149]), .B(
        b11_OFWNT9L_8tZ[5]), .C(b4_nUAi[448]), .D(b4_nUAi[447]), .Y(
        b3_P_F_6_am_62));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[149]), .B(
        b11_OFWNT9L_8tZ[5]), .C(b4_nUAi[447]), .D(b4_nUAi[448]), .Y(
        b3_P_F_6_bm_62));
    
endmodule


module b8_1LbcQDr1_x_63_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [91:91] mdiclink_reg;
input  [63:63] b11_OFWNT9L_8tZ;
input  [275:273] b4_nUAi;
output [91:91] b6_2ZTGIf;

    wire b3_P_F_6_bm_23, b3_P_F_6_am_23, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_23), .B(
        b4_nUAi[275]), .C(b3_P_F_6_am_23), .Y(b6_2ZTGIf[91]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[91]), .B(
        b11_OFWNT9L_8tZ[63]), .C(b4_nUAi[274]), .D(b4_nUAi[273]), .Y(
        b3_P_F_6_am_23));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[91]), .B(
        b11_OFWNT9L_8tZ[63]), .C(b4_nUAi[273]), .D(b4_nUAi[274]), .Y(
        b3_P_F_6_bm_23));
    
endmodule


module b8_1LbcQDr1_x_149_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [5:5] mdiclink_reg;
input  [149:149] b11_OFWNT9L_8tZ;
input  [17:15] b4_nUAi;
output [5:5] b6_2ZTGIf;

    wire b3_P_F_6_bm_74, b3_P_F_6_am_74, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_74), .B(
        b4_nUAi[17]), .C(b3_P_F_6_am_74), .Y(b6_2ZTGIf[5]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[5]), .B(
        b11_OFWNT9L_8tZ[149]), .C(b4_nUAi[16]), .D(b4_nUAi[15]), .Y(
        b3_P_F_6_am_74));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[5]), .B(
        b11_OFWNT9L_8tZ[149]), .C(b4_nUAi[15]), .D(b4_nUAi[16]), .Y(
        b3_P_F_6_bm_74));
    
endmodule


module b8_1LbcQDr1_x_6_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [148:148] mdiclink_reg;
input  [6:6] b11_OFWNT9L_8tZ;
input  [445:444] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[148]), .B(
        b11_OFWNT9L_8tZ[6]), .C(b4_nUAi[445]), .D(b4_nUAi[444]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[148]), .B(
        b11_OFWNT9L_8tZ[6]), .C(b4_nUAi[445]), .D(b4_nUAi[444]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_64_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [90:90] mdiclink_reg;
input  [64:64] b11_OFWNT9L_8tZ;
input  [271:270] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[90]), .B(
        b11_OFWNT9L_8tZ[64]), .C(b4_nUAi[271]), .D(b4_nUAi[270]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[90]), .B(
        b11_OFWNT9L_8tZ[64]), .C(b4_nUAi[271]), .D(b4_nUAi[270]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_22_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [132:132] mdiclink_reg;
input  [22:22] b11_OFWNT9L_8tZ;
input  [398:396] b4_nUAi;
output [132:132] b6_2ZTGIf;

    wire b3_P_F_6_bm_58, b3_P_F_6_am_58, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_58), .B(
        b4_nUAi[398]), .C(b3_P_F_6_am_58), .Y(b6_2ZTGIf[132]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[132]), .B(
        b11_OFWNT9L_8tZ[22]), .C(b4_nUAi[397]), .D(b4_nUAi[396]), .Y(
        b3_P_F_6_am_58));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[132]), .B(
        b11_OFWNT9L_8tZ[22]), .C(b4_nUAi[396]), .D(b4_nUAi[397]), .Y(
        b3_P_F_6_bm_58));
    
endmodule


module b8_1LbcQDr1_x_7_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [147:147] mdiclink_reg;
input  [7:7] b11_OFWNT9L_8tZ;
input  [443:441] b4_nUAi;
output [147:147] b6_2ZTGIf;

    wire b3_P_F_6_bm_63, b3_P_F_6_am_63, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_63), .B(
        b4_nUAi[443]), .C(b3_P_F_6_am_63), .Y(b6_2ZTGIf[147]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[147]), .B(
        b11_OFWNT9L_8tZ[7]), .C(b4_nUAi[442]), .D(b4_nUAi[441]), .Y(
        b3_P_F_6_am_63));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[147]), .B(
        b11_OFWNT9L_8tZ[7]), .C(b4_nUAi[441]), .D(b4_nUAi[442]), .Y(
        b3_P_F_6_bm_63));
    
endmodule


module b8_1LbcQDr1_x_77_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [77:77] mdiclink_reg;
input  [77:77] b11_OFWNT9L_8tZ;
input  [233:231] b4_nUAi;
output [77:77] b6_2ZTGIf;

    wire b3_P_F_6_bm_11, b3_P_F_6_am_11, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_11), .B(
        b4_nUAi[233]), .C(b3_P_F_6_am_11), .Y(b6_2ZTGIf[77]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[77]), .B(
        b11_OFWNT9L_8tZ[77]), .C(b4_nUAi[232]), .D(b4_nUAi[231]), .Y(
        b3_P_F_6_am_11));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[77]), .B(
        b11_OFWNT9L_8tZ[77]), .C(b4_nUAi[231]), .D(b4_nUAi[232]), .Y(
        b3_P_F_6_bm_11));
    
endmodule


module b8_1LbcQDr1_x_137_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [17:17] mdiclink_reg;
input  [137:137] b11_OFWNT9L_8tZ;
input  [52:51] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[17]), .B(
        b11_OFWNT9L_8tZ[137]), .C(b4_nUAi[52]), .D(b4_nUAi[51]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[17]), .B(
        b11_OFWNT9L_8tZ[137]), .C(b4_nUAi[52]), .D(b4_nUAi[51]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_100_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [54:54] mdiclink_reg;
input  [100:100] b11_OFWNT9L_8tZ;
input  [164:162] b4_nUAi;
output [54:54] b6_2ZTGIf;

    wire b3_P_F_6_bm_6, b3_P_F_6_am_6, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_6), .B(
        b4_nUAi[164]), .C(b3_P_F_6_am_6), .Y(b6_2ZTGIf[54]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[54]), .B(
        b11_OFWNT9L_8tZ[100]), .C(b4_nUAi[163]), .D(b4_nUAi[162]), .Y(
        b3_P_F_6_am_6));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[54]), .B(
        b11_OFWNT9L_8tZ[100]), .C(b4_nUAi[162]), .D(b4_nUAi[163]), .Y(
        b3_P_F_6_bm_6));
    
endmodule


module b8_1LbcQDr1_x_152_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [2:2] mdiclink_reg;
input  [152:152] b11_OFWNT9L_8tZ;
input  [7:6] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[2]), .B(
        b11_OFWNT9L_8tZ[152]), .C(b4_nUAi[7]), .D(b4_nUAi[6]), .Y(N_27)
        );
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[2]), .B(
        b11_OFWNT9L_8tZ[152]), .C(b4_nUAi[7]), .D(b4_nUAi[6]), .Y(N_25)
        );
    
endmodule


module b8_1LbcQDr1_x_97_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [57:57] mdiclink_reg;
input  [97:97] b11_OFWNT9L_8tZ;
input  [173:171] b4_nUAi;
output [57:57] b6_2ZTGIf;

    wire b3_P_F_6_bm_4, b3_P_F_6_am_4, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_4), .B(
        b4_nUAi[173]), .C(b3_P_F_6_am_4), .Y(b6_2ZTGIf[57]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[57]), .B(
        b11_OFWNT9L_8tZ[97]), .C(b4_nUAi[172]), .D(b4_nUAi[171]), .Y(
        b3_P_F_6_am_4));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[57]), .B(
        b11_OFWNT9L_8tZ[97]), .C(b4_nUAi[171]), .D(b4_nUAi[172]), .Y(
        b3_P_F_6_bm_4));
    
endmodule


module b8_1LbcQDr1_x_14_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [140:140] mdiclink_reg;
input  [14:14] b11_OFWNT9L_8tZ;
input  [422:420] b4_nUAi;
output [140:140] b6_2ZTGIf;

    wire b3_P_F_6_bm_52, b3_P_F_6_am_52, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_52), .B(
        b4_nUAi[422]), .C(b3_P_F_6_am_52), .Y(b6_2ZTGIf[140]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[140]), .B(
        b11_OFWNT9L_8tZ[14]), .C(b4_nUAi[421]), .D(b4_nUAi[420]), .Y(
        b3_P_F_6_am_52));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[140]), .B(
        b11_OFWNT9L_8tZ[14]), .C(b4_nUAi[420]), .D(b4_nUAi[421]), .Y(
        b3_P_F_6_bm_52));
    
endmodule


module b8_1LbcQDr1_x_116_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [38:38] mdiclink_reg;
input  [116:116] b11_OFWNT9L_8tZ;
input  [116:114] b4_nUAi;
output [38:38] b6_2ZTGIf;

    wire b3_P_F_6_bm_93, b3_P_F_6_am_93, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_93), .B(
        b4_nUAi[116]), .C(b3_P_F_6_am_93), .Y(b6_2ZTGIf[38]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[38]), .B(
        b11_OFWNT9L_8tZ[116]), .C(b4_nUAi[115]), .D(b4_nUAi[114]), .Y(
        b3_P_F_6_am_93));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[38]), .B(
        b11_OFWNT9L_8tZ[116]), .C(b4_nUAi[114]), .D(b4_nUAi[115]), .Y(
        b3_P_F_6_bm_93));
    
endmodule


module b8_1LbcQDr1_x_68_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [86:86] mdiclink_reg;
input  [68:68] b11_OFWNT9L_8tZ;
input  [260:258] b4_nUAi;
output [86:86] b6_2ZTGIf;

    wire b3_P_F_6_bm_26, b3_P_F_6_am_26, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_26), .B(
        b4_nUAi[260]), .C(b3_P_F_6_am_26), .Y(b6_2ZTGIf[86]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[86]), .B(
        b11_OFWNT9L_8tZ[68]), .C(b4_nUAi[259]), .D(b4_nUAi[258]), .Y(
        b3_P_F_6_am_26));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[86]), .B(
        b11_OFWNT9L_8tZ[68]), .C(b4_nUAi[258]), .D(b4_nUAi[259]), .Y(
        b3_P_F_6_bm_26));
    
endmodule


module b8_1LbcQDr1_x_112_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [42:42] mdiclink_reg;
input  [112:112] b11_OFWNT9L_8tZ;
input  [127:126] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[42]), .B(
        b11_OFWNT9L_8tZ[112]), .C(b4_nUAi[127]), .D(b4_nUAi[126]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[42]), .B(
        b11_OFWNT9L_8tZ[112]), .C(b4_nUAi[127]), .D(b4_nUAi[126]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_19_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [135:135] mdiclink_reg;
input  [19:19] b11_OFWNT9L_8tZ;
input  [407:405] b4_nUAi;
output [135:135] b6_2ZTGIf;

    wire b3_P_F_6_bm_55, b3_P_F_6_am_55, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_55), .B(
        b4_nUAi[407]), .C(b3_P_F_6_am_55), .Y(b6_2ZTGIf[135]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[135]), .B(
        b11_OFWNT9L_8tZ[19]), .C(b4_nUAi[406]), .D(b4_nUAi[405]), .Y(
        b3_P_F_6_am_55));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[135]), .B(
        b11_OFWNT9L_8tZ[19]), .C(b4_nUAi[405]), .D(b4_nUAi[406]), .Y(
        b3_P_F_6_bm_55));
    
endmodule


module b8_1LbcQDr1_x_115_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [39:39] mdiclink_reg;
input  [115:115] b11_OFWNT9L_8tZ;
input  [119:117] b4_nUAi;
output [39:39] b6_2ZTGIf;

    wire b3_P_F_6_bm_92, b3_P_F_6_am_92, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_92), .B(
        b4_nUAi[119]), .C(b3_P_F_6_am_92), .Y(b6_2ZTGIf[39]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[39]), .B(
        b11_OFWNT9L_8tZ[115]), .C(b4_nUAi[118]), .D(b4_nUAi[117]), .Y(
        b3_P_F_6_am_92));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[39]), .B(
        b11_OFWNT9L_8tZ[115]), .C(b4_nUAi[117]), .D(b4_nUAi[118]), .Y(
        b3_P_F_6_bm_92));
    
endmodule


module b8_1LbcQDr1_x_13_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [141:141] mdiclink_reg;
input  [13:13] b11_OFWNT9L_8tZ;
input  [425:423] b4_nUAi;
output [141:141] b6_2ZTGIf;

    wire b3_P_F_6_bm_51, b3_P_F_6_am_51, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_51), .B(
        b4_nUAi[425]), .C(b3_P_F_6_am_51), .Y(b6_2ZTGIf[141]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[141]), .B(
        b11_OFWNT9L_8tZ[13]), .C(b4_nUAi[424]), .D(b4_nUAi[423]), .Y(
        b3_P_F_6_am_51));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[141]), .B(
        b11_OFWNT9L_8tZ[13]), .C(b4_nUAi[423]), .D(b4_nUAi[424]), .Y(
        b3_P_F_6_bm_51));
    
endmodule


module b8_1LbcQDr1_x_15_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [139:139] mdiclink_reg;
input  [15:15] b11_OFWNT9L_8tZ;
input  [419:417] b4_nUAi;
output [139:139] b6_2ZTGIf;

    wire b3_P_F_6_bm_53, b3_P_F_6_am_53, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_53), .B(
        b4_nUAi[419]), .C(b3_P_F_6_am_53), .Y(b6_2ZTGIf[139]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[139]), .B(
        b11_OFWNT9L_8tZ[15]), .C(b4_nUAi[418]), .D(b4_nUAi[417]), .Y(
        b3_P_F_6_am_53));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[139]), .B(
        b11_OFWNT9L_8tZ[15]), .C(b4_nUAi[417]), .D(b4_nUAi[418]), .Y(
        b3_P_F_6_bm_53));
    
endmodule


module b8_1LbcQDr1_x_42_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [112:112] mdiclink_reg;
input  [42:42] b11_OFWNT9L_8tZ;
input  [337:336] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[112]), .B(
        b11_OFWNT9L_8tZ[42]), .C(b4_nUAi[337]), .D(b4_nUAi[336]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[112]), .B(
        b11_OFWNT9L_8tZ[42]), .C(b4_nUAi[337]), .D(b4_nUAi[336]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_0_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf,
       b7_PSyi3wy
    );
input  [154:154] mdiclink_reg;
input  [0:0] b11_OFWNT9L_8tZ;
input  [463:462] b4_nUAi;
output [154:154] b6_2ZTGIf;
input  b7_PSyi3wy;

    wire b3_P_F_6_bm_59, b3_P_F_6_am_59, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_59), .B(
        b7_PSyi3wy), .C(b3_P_F_6_am_59), .Y(b6_2ZTGIf[154]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[154]), .B(
        b11_OFWNT9L_8tZ[0]), .C(b4_nUAi[463]), .D(b4_nUAi[462]), .Y(
        b3_P_F_6_am_59));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[154]), .B(
        b11_OFWNT9L_8tZ[0]), .C(b4_nUAi[462]), .D(b4_nUAi[463]), .Y(
        b3_P_F_6_bm_59));
    
endmodule


module b8_1LbcQDr1_x_52_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [102:102] mdiclink_reg;
input  [52:52] b11_OFWNT9L_8tZ;
input  [308:306] b4_nUAi;
output [102:102] b6_2ZTGIf;

    wire b3_P_F_6_bm_36, b3_P_F_6_am_36, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_36), .B(
        b4_nUAi[308]), .C(b3_P_F_6_am_36), .Y(b6_2ZTGIf[102]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[102]), .B(
        b11_OFWNT9L_8tZ[52]), .C(b4_nUAi[307]), .D(b4_nUAi[306]), .Y(
        b3_P_F_6_am_36));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[102]), .B(
        b11_OFWNT9L_8tZ[52]), .C(b4_nUAi[306]), .D(b4_nUAi[307]), .Y(
        b3_P_F_6_bm_36));
    
endmodule


module b8_1LbcQDr1_x_16_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [138:138] mdiclink_reg;
input  [16:16] b11_OFWNT9L_8tZ;
input  [415:414] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[138]), .B(
        b11_OFWNT9L_8tZ[16]), .C(b4_nUAi[415]), .D(b4_nUAi[414]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[138]), .B(
        b11_OFWNT9L_8tZ[16]), .C(b4_nUAi[415]), .D(b4_nUAi[414]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_17_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [137:137] mdiclink_reg;
input  [17:17] b11_OFWNT9L_8tZ;
input  [413:411] b4_nUAi;
output [137:137] b6_2ZTGIf;

    wire b3_P_F_6_bm_54, b3_P_F_6_am_54, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_54), .B(
        b4_nUAi[413]), .C(b3_P_F_6_am_54), .Y(b6_2ZTGIf[137]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[137]), .B(
        b11_OFWNT9L_8tZ[17]), .C(b4_nUAi[412]), .D(b4_nUAi[411]), .Y(
        b3_P_F_6_am_54));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[137]), .B(
        b11_OFWNT9L_8tZ[17]), .C(b4_nUAi[411]), .D(b4_nUAi[412]), .Y(
        b3_P_F_6_bm_54));
    
endmodule


module b8_1LbcQDr1_x_128_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [26:26] mdiclink_reg;
input  [128:128] b11_OFWNT9L_8tZ;
input  [79:78] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[26]), .B(
        b11_OFWNT9L_8tZ[128]), .C(b4_nUAi[79]), .D(b4_nUAi[78]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[26]), .B(
        b11_OFWNT9L_8tZ[128]), .C(b4_nUAi[79]), .D(b4_nUAi[78]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_154_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [0:0] mdiclink_reg;
input  [154:154] b11_OFWNT9L_8tZ;
input  [1:0] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[0]), .B(
        b11_OFWNT9L_8tZ[154]), .C(b4_nUAi[1]), .D(b4_nUAi[0]), .Y(N_27)
        );
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[0]), .B(
        b11_OFWNT9L_8tZ[154]), .C(b4_nUAi[1]), .D(b4_nUAi[0]), .Y(N_25)
        );
    
endmodule


module b8_1LbcQDr1_x_24_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [130:130] mdiclink_reg;
input  [24:24] b11_OFWNT9L_8tZ;
input  [391:390] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[130]), .B(
        b11_OFWNT9L_8tZ[24]), .C(b4_nUAi[391]), .D(b4_nUAi[390]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[130]), .B(
        b11_OFWNT9L_8tZ[24]), .C(b4_nUAi[391]), .D(b4_nUAi[390]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_88_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [66:66] mdiclink_reg;
input  [88:88] b11_OFWNT9L_8tZ;
input  [199:198] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[66]), .B(
        b11_OFWNT9L_8tZ[88]), .C(b4_nUAi[199]), .D(b4_nUAi[198]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[66]), .B(
        b11_OFWNT9L_8tZ[88]), .C(b4_nUAi[199]), .D(b4_nUAi[198]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_39_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [115:115] mdiclink_reg;
input  [39:39] b11_OFWNT9L_8tZ;
input  [346:345] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[115]), .B(
        b11_OFWNT9L_8tZ[39]), .C(b4_nUAi[346]), .D(b4_nUAi[345]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[115]), .B(
        b11_OFWNT9L_8tZ[39]), .C(b4_nUAi[346]), .D(b4_nUAi[345]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_49_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [105:105] mdiclink_reg;
input  [49:49] b11_OFWNT9L_8tZ;
input  [317:315] b4_nUAi;
output [105:105] b6_2ZTGIf;

    wire b3_P_F_6_bm_34, b3_P_F_6_am_34, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_34), .B(
        b4_nUAi[317]), .C(b3_P_F_6_am_34), .Y(b6_2ZTGIf[105]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[105]), .B(
        b11_OFWNT9L_8tZ[49]), .C(b4_nUAi[316]), .D(b4_nUAi[315]), .Y(
        b3_P_F_6_am_34));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[105]), .B(
        b11_OFWNT9L_8tZ[49]), .C(b4_nUAi[315]), .D(b4_nUAi[316]), .Y(
        b3_P_F_6_bm_34));
    
endmodule


module b8_1LbcQDr1_x_56_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [98:98] mdiclink_reg;
input  [56:56] b11_OFWNT9L_8tZ;
input  [295:294] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[98]), .B(
        b11_OFWNT9L_8tZ[56]), .C(b4_nUAi[295]), .D(b4_nUAi[294]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[98]), .B(
        b11_OFWNT9L_8tZ[56]), .C(b4_nUAi[295]), .D(b4_nUAi[294]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_71_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [83:83] mdiclink_reg;
input  [71:71] b11_OFWNT9L_8tZ;
input  [250:249] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[83]), .B(
        b11_OFWNT9L_8tZ[71]), .C(b4_nUAi[250]), .D(b4_nUAi[249]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[83]), .B(
        b11_OFWNT9L_8tZ[71]), .C(b4_nUAi[250]), .D(b4_nUAi[249]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_30_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [124:124] mdiclink_reg;
input  [30:30] b11_OFWNT9L_8tZ;
input  [374:372] b4_nUAi;
output [124:124] b6_2ZTGIf;

    wire b3_P_F_6_bm_42, b3_P_F_6_am_42, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_42), .B(
        b4_nUAi[374]), .C(b3_P_F_6_am_42), .Y(b6_2ZTGIf[124]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[124]), .B(
        b11_OFWNT9L_8tZ[30]), .C(b4_nUAi[373]), .D(b4_nUAi[372]), .Y(
        b3_P_F_6_am_42));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[124]), .B(
        b11_OFWNT9L_8tZ[30]), .C(b4_nUAi[372]), .D(b4_nUAi[373]), .Y(
        b3_P_F_6_bm_42));
    
endmodule


module b8_1LbcQDr1_x_107_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [47:47] mdiclink_reg;
input  [107:107] b11_OFWNT9L_8tZ;
input  [143:141] b4_nUAi;
output [47:47] b6_2ZTGIf;

    wire b3_P_F_6_bm_86, b3_P_F_6_am_86, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_86), .B(
        b4_nUAi[143]), .C(b3_P_F_6_am_86), .Y(b6_2ZTGIf[47]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[47]), .B(
        b11_OFWNT9L_8tZ[107]), .C(b4_nUAi[142]), .D(b4_nUAi[141]), .Y(
        b3_P_F_6_am_86));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[47]), .B(
        b11_OFWNT9L_8tZ[107]), .C(b4_nUAi[141]), .D(b4_nUAi[142]), .Y(
        b3_P_F_6_bm_86));
    
endmodule


module b8_1LbcQDr1_x_35_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [119:119] mdiclink_reg;
input  [35:35] b11_OFWNT9L_8tZ;
input  [359:357] b4_nUAi;
output [119:119] b6_2ZTGIf;

    wire b3_P_F_6_bm_45, b3_P_F_6_am_45, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_45), .B(
        b4_nUAi[359]), .C(b3_P_F_6_am_45), .Y(b6_2ZTGIf[119]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[119]), .B(
        b11_OFWNT9L_8tZ[35]), .C(b4_nUAi[358]), .D(b4_nUAi[357]), .Y(
        b3_P_F_6_am_45));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[119]), .B(
        b11_OFWNT9L_8tZ[35]), .C(b4_nUAi[357]), .D(b4_nUAi[358]), .Y(
        b3_P_F_6_bm_45));
    
endmodule


module b8_1LbcQDr1_x_28_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [126:126] mdiclink_reg;
input  [28:28] b11_OFWNT9L_8tZ;
input  [380:378] b4_nUAi;
output [126:126] b6_2ZTGIf;

    wire b3_P_F_6_bm_40, b3_P_F_6_am_40, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_40), .B(
        b4_nUAi[380]), .C(b3_P_F_6_am_40), .Y(b6_2ZTGIf[126]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[126]), .B(
        b11_OFWNT9L_8tZ[28]), .C(b4_nUAi[379]), .D(b4_nUAi[378]), .Y(
        b3_P_F_6_am_40));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[126]), .B(
        b11_OFWNT9L_8tZ[28]), .C(b4_nUAi[378]), .D(b4_nUAi[379]), .Y(
        b3_P_F_6_bm_40));
    
endmodule


module b8_1LbcQDr1_x_23_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [131:131] mdiclink_reg;
input  [23:23] b11_OFWNT9L_8tZ;
input  [394:393] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[131]), .B(
        b11_OFWNT9L_8tZ[23]), .C(b4_nUAi[394]), .D(b4_nUAi[393]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[131]), .B(
        b11_OFWNT9L_8tZ[23]), .C(b4_nUAi[394]), .D(b4_nUAi[393]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_45_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [109:109] mdiclink_reg;
input  [45:45] b11_OFWNT9L_8tZ;
input  [329:327] b4_nUAi;
output [109:109] b6_2ZTGIf;

    wire b3_P_F_6_bm_31, b3_P_F_6_am_31, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_31), .B(
        b4_nUAi[329]), .C(b3_P_F_6_am_31), .Y(b6_2ZTGIf[109]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[109]), .B(
        b11_OFWNT9L_8tZ[45]), .C(b4_nUAi[328]), .D(b4_nUAi[327]), .Y(
        b3_P_F_6_am_31));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[109]), .B(
        b11_OFWNT9L_8tZ[45]), .C(b4_nUAi[327]), .D(b4_nUAi[328]), .Y(
        b3_P_F_6_bm_31));
    
endmodule


module b8_1LbcQDr1_x_36_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [118:118] mdiclink_reg;
input  [36:36] b11_OFWNT9L_8tZ;
input  [356:354] b4_nUAi;
output [118:118] b6_2ZTGIf;

    wire b3_P_F_6_bm_46, b3_P_F_6_am_46, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_46), .B(
        b4_nUAi[356]), .C(b3_P_F_6_am_46), .Y(b6_2ZTGIf[118]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[118]), .B(
        b11_OFWNT9L_8tZ[36]), .C(b4_nUAi[355]), .D(b4_nUAi[354]), .Y(
        b3_P_F_6_am_46));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[118]), .B(
        b11_OFWNT9L_8tZ[36]), .C(b4_nUAi[354]), .D(b4_nUAi[355]), .Y(
        b3_P_F_6_bm_46));
    
endmodule


module b8_1LbcQDr1_x_55_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [99:99] mdiclink_reg;
input  [55:55] b11_OFWNT9L_8tZ;
input  [298:297] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[99]), .B(
        b11_OFWNT9L_8tZ[55]), .C(b4_nUAi[298]), .D(b4_nUAi[297]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[99]), .B(
        b11_OFWNT9L_8tZ[55]), .C(b4_nUAi[298]), .D(b4_nUAi[297]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_119_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [35:35] mdiclink_reg;
input  [119:119] b11_OFWNT9L_8tZ;
input  [106:105] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[35]), .B(
        b11_OFWNT9L_8tZ[119]), .C(b4_nUAi[106]), .D(b4_nUAi[105]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[35]), .B(
        b11_OFWNT9L_8tZ[119]), .C(b4_nUAi[106]), .D(b4_nUAi[105]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_46_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [108:108] mdiclink_reg;
input  [46:46] b11_OFWNT9L_8tZ;
input  [326:324] b4_nUAi;
output [108:108] b6_2ZTGIf;

    wire b3_P_F_6_bm_32, b3_P_F_6_am_32, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_32), .B(
        b4_nUAi[326]), .C(b3_P_F_6_am_32), .Y(b6_2ZTGIf[108]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[108]), .B(
        b11_OFWNT9L_8tZ[46]), .C(b4_nUAi[325]), .D(b4_nUAi[324]), .Y(
        b3_P_F_6_am_32));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[108]), .B(
        b11_OFWNT9L_8tZ[46]), .C(b4_nUAi[324]), .D(b4_nUAi[325]), .Y(
        b3_P_F_6_bm_32));
    
endmodule


module b8_1LbcQDr1_x_151_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [3:3] mdiclink_reg;
input  [151:151] b11_OFWNT9L_8tZ;
input  [10:9] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[3]), .B(
        b11_OFWNT9L_8tZ[151]), .C(b4_nUAi[10]), .D(b4_nUAi[9]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[3]), .B(
        b11_OFWNT9L_8tZ[151]), .C(b4_nUAi[10]), .D(b4_nUAi[9]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_37_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [117:117] mdiclink_reg;
input  [37:37] b11_OFWNT9L_8tZ;
input  [353:351] b4_nUAi;
output [117:117] b6_2ZTGIf;

    wire b3_P_F_6_bm_47, b3_P_F_6_am_47, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_47), .B(
        b4_nUAi[353]), .C(b3_P_F_6_am_47), .Y(b6_2ZTGIf[117]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[117]), .B(
        b11_OFWNT9L_8tZ[37]), .C(b4_nUAi[352]), .D(b4_nUAi[351]), .Y(
        b3_P_F_6_am_47));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[117]), .B(
        b11_OFWNT9L_8tZ[37]), .C(b4_nUAi[351]), .D(b4_nUAi[352]), .Y(
        b3_P_F_6_bm_47));
    
endmodule


module b8_1LbcQDr1_x_11_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [143:143] mdiclink_reg;
input  [11:11] b11_OFWNT9L_8tZ;
input  [431:429] b4_nUAi;
output [143:143] b6_2ZTGIf;

    wire b3_P_F_6_bm_49, b3_P_F_6_am_49, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_49), .B(
        b4_nUAi[431]), .C(b3_P_F_6_am_49), .Y(b6_2ZTGIf[143]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[143]), .B(
        b11_OFWNT9L_8tZ[11]), .C(b4_nUAi[430]), .D(b4_nUAi[429]), .Y(
        b3_P_F_6_am_49));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[143]), .B(
        b11_OFWNT9L_8tZ[11]), .C(b4_nUAi[429]), .D(b4_nUAi[430]), .Y(
        b3_P_F_6_bm_49));
    
endmodule


module b8_1LbcQDr1_x_47_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [107:107] mdiclink_reg;
input  [47:47] b11_OFWNT9L_8tZ;
input  [323:321] b4_nUAi;
output [107:107] b6_2ZTGIf;

    wire b3_P_F_6_bm_33, b3_P_F_6_am_33, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_33), .B(
        b4_nUAi[323]), .C(b3_P_F_6_am_33), .Y(b6_2ZTGIf[107]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[107]), .B(
        b11_OFWNT9L_8tZ[47]), .C(b4_nUAi[322]), .D(b4_nUAi[321]), .Y(
        b3_P_F_6_am_33));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[107]), .B(
        b11_OFWNT9L_8tZ[47]), .C(b4_nUAi[321]), .D(b4_nUAi[322]), .Y(
        b3_P_F_6_bm_33));
    
endmodule


module b8_1LbcQDr1_x_44_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [110:110] mdiclink_reg;
input  [44:44] b11_OFWNT9L_8tZ;
input  [332:330] b4_nUAi;
output [110:110] b6_2ZTGIf;

    wire b3_P_F_6_bm_30, b3_P_F_6_am_30, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_30), .B(
        b4_nUAi[332]), .C(b3_P_F_6_am_30), .Y(b6_2ZTGIf[110]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[110]), .B(
        b11_OFWNT9L_8tZ[44]), .C(b4_nUAi[331]), .D(b4_nUAi[330]), .Y(
        b3_P_F_6_am_30));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[110]), .B(
        b11_OFWNT9L_8tZ[44]), .C(b4_nUAi[330]), .D(b4_nUAi[331]), .Y(
        b3_P_F_6_bm_30));
    
endmodule


module b8_1LbcQDr1_x_54_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [100:100] mdiclink_reg;
input  [54:54] b11_OFWNT9L_8tZ;
input  [302:300] b4_nUAi;
output [100:100] b6_2ZTGIf;

    wire b3_P_F_6_bm_38, b3_P_F_6_am_38, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_38), .B(
        b4_nUAi[302]), .C(b3_P_F_6_am_38), .Y(b6_2ZTGIf[100]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[100]), .B(
        b11_OFWNT9L_8tZ[54]), .C(b4_nUAi[301]), .D(b4_nUAi[300]), .Y(
        b3_P_F_6_am_38));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[100]), .B(
        b11_OFWNT9L_8tZ[54]), .C(b4_nUAi[300]), .D(b4_nUAi[301]), .Y(
        b3_P_F_6_bm_38));
    
endmodule


module b8_1LbcQDr1_x_73_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [81:81] mdiclink_reg;
input  [73:73] b11_OFWNT9L_8tZ;
input  [244:243] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[81]), .B(
        b11_OFWNT9L_8tZ[73]), .C(b4_nUAi[244]), .D(b4_nUAi[243]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[81]), .B(
        b11_OFWNT9L_8tZ[73]), .C(b4_nUAi[244]), .D(b4_nUAi[243]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_74_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [80:80] mdiclink_reg;
input  [74:74] b11_OFWNT9L_8tZ;
input  [241:240] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[80]), .B(
        b11_OFWNT9L_8tZ[74]), .C(b4_nUAi[241]), .D(b4_nUAi[240]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[80]), .B(
        b11_OFWNT9L_8tZ[74]), .C(b4_nUAi[241]), .D(b4_nUAi[240]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_122_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [32:32] mdiclink_reg;
input  [122:122] b11_OFWNT9L_8tZ;
input  [97:96] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[32]), .B(
        b11_OFWNT9L_8tZ[122]), .C(b4_nUAi[97]), .D(b4_nUAi[96]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[32]), .B(
        b11_OFWNT9L_8tZ[122]), .C(b4_nUAi[97]), .D(b4_nUAi[96]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_43_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [111:111] mdiclink_reg;
input  [43:43] b11_OFWNT9L_8tZ;
input  [335:333] b4_nUAi;
output [111:111] b6_2ZTGIf;

    wire b3_P_F_6_bm_29, b3_P_F_6_am_29, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_29), .B(
        b4_nUAi[335]), .C(b3_P_F_6_am_29), .Y(b6_2ZTGIf[111]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[111]), .B(
        b11_OFWNT9L_8tZ[43]), .C(b4_nUAi[334]), .D(b4_nUAi[333]), .Y(
        b3_P_F_6_am_29));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[111]), .B(
        b11_OFWNT9L_8tZ[43]), .C(b4_nUAi[333]), .D(b4_nUAi[334]), .Y(
        b3_P_F_6_bm_29));
    
endmodule


module b8_1LbcQDr1_x_131_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [23:23] mdiclink_reg;
input  [131:131] b11_OFWNT9L_8tZ;
input  [71:69] b4_nUAi;
output [23:23] b6_2ZTGIf;

    wire b3_P_F_6_bm_82, b3_P_F_6_am_82, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_82), .B(
        b4_nUAi[71]), .C(b3_P_F_6_am_82), .Y(b6_2ZTGIf[23]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[23]), .B(
        b11_OFWNT9L_8tZ[131]), .C(b4_nUAi[70]), .D(b4_nUAi[69]), .Y(
        b3_P_F_6_am_82));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[23]), .B(
        b11_OFWNT9L_8tZ[131]), .C(b4_nUAi[69]), .D(b4_nUAi[70]), .Y(
        b3_P_F_6_bm_82));
    
endmodule


module b8_1LbcQDr1_x_91_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [63:63] mdiclink_reg;
input  [91:91] b11_OFWNT9L_8tZ;
input  [191:189] b4_nUAi;
output [63:63] b6_2ZTGIf;

    wire b3_P_F_6_bm_net_1, b3_P_F_6_am_net_1, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_net_1), .B(
        b4_nUAi[191]), .C(b3_P_F_6_am_net_1), .Y(b6_2ZTGIf[63]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[63]), .B(
        b11_OFWNT9L_8tZ[91]), .C(b4_nUAi[190]), .D(b4_nUAi[189]), .Y(
        b3_P_F_6_am_net_1));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[63]), .B(
        b11_OFWNT9L_8tZ[91]), .C(b4_nUAi[189]), .D(b4_nUAi[190]), .Y(
        b3_P_F_6_bm_net_1));
    
endmodule


module b8_1LbcQDr1_x_53_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [101:101] mdiclink_reg;
input  [53:53] b11_OFWNT9L_8tZ;
input  [305:303] b4_nUAi;
output [101:101] b6_2ZTGIf;

    wire b3_P_F_6_bm_37, b3_P_F_6_am_37, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_37), .B(
        b4_nUAi[305]), .C(b3_P_F_6_am_37), .Y(b6_2ZTGIf[101]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[101]), .B(
        b11_OFWNT9L_8tZ[53]), .C(b4_nUAi[304]), .D(b4_nUAi[303]), .Y(
        b3_P_F_6_am_37));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[101]), .B(
        b11_OFWNT9L_8tZ[53]), .C(b4_nUAi[303]), .D(b4_nUAi[304]), .Y(
        b3_P_F_6_bm_37));
    
endmodule


module b8_1LbcQDr1_x_21_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [133:133] mdiclink_reg;
input  [21:21] b11_OFWNT9L_8tZ;
input  [401:399] b4_nUAi;
output [133:133] b6_2ZTGIf;

    wire b3_P_F_6_bm_57, b3_P_F_6_am_57, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_57), .B(
        b4_nUAi[401]), .C(b3_P_F_6_am_57), .Y(b6_2ZTGIf[133]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[133]), .B(
        b11_OFWNT9L_8tZ[21]), .C(b4_nUAi[400]), .D(b4_nUAi[399]), .Y(
        b3_P_F_6_am_57));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[133]), .B(
        b11_OFWNT9L_8tZ[21]), .C(b4_nUAi[399]), .D(b4_nUAi[400]), .Y(
        b3_P_F_6_bm_57));
    
endmodule


module b8_1LbcQDr1_x_59_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [95:95] mdiclink_reg;
input  [59:59] b11_OFWNT9L_8tZ;
input  [287:285] b4_nUAi;
output [95:95] b6_2ZTGIf;

    wire b3_P_F_6_bm_19, b3_P_F_6_am_19, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_19), .B(
        b4_nUAi[287]), .C(b3_P_F_6_am_19), .Y(b6_2ZTGIf[95]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[95]), .B(
        b11_OFWNT9L_8tZ[59]), .C(b4_nUAi[286]), .D(b4_nUAi[285]), .Y(
        b3_P_F_6_am_19));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[95]), .B(
        b11_OFWNT9L_8tZ[59]), .C(b4_nUAi[285]), .D(b4_nUAi[286]), .Y(
        b3_P_F_6_bm_19));
    
endmodule


module b8_1LbcQDr1_x_146_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [8:8] mdiclink_reg;
input  [146:146] b11_OFWNT9L_8tZ;
input  [25:24] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[8]), .B(
        b11_OFWNT9L_8tZ[146]), .C(b4_nUAi[25]), .D(b4_nUAi[24]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[8]), .B(
        b11_OFWNT9L_8tZ[146]), .C(b4_nUAi[25]), .D(b4_nUAi[24]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_133_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [21:21] mdiclink_reg;
input  [133:133] b11_OFWNT9L_8tZ;
input  [65:63] b4_nUAi;
output [21:21] b6_2ZTGIf;

    wire b3_P_F_6_bm_84, b3_P_F_6_am_84, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_84), .B(
        b4_nUAi[65]), .C(b3_P_F_6_am_84), .Y(b6_2ZTGIf[21]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[21]), .B(
        b11_OFWNT9L_8tZ[133]), .C(b4_nUAi[64]), .D(b4_nUAi[63]), .Y(
        b3_P_F_6_am_84));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[21]), .B(
        b11_OFWNT9L_8tZ[133]), .C(b4_nUAi[63]), .D(b4_nUAi[64]), .Y(
        b3_P_F_6_bm_84));
    
endmodule


module b8_1LbcQDr1_x_93_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [61:61] mdiclink_reg;
input  [93:93] b11_OFWNT9L_8tZ;
input  [185:183] b4_nUAi;
output [61:61] b6_2ZTGIf;

    wire b3_P_F_6_bm_1, b3_P_F_6_am_1, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_1), .B(
        b4_nUAi[185]), .C(b3_P_F_6_am_1), .Y(b6_2ZTGIf[61]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[61]), .B(
        b11_OFWNT9L_8tZ[93]), .C(b4_nUAi[184]), .D(b4_nUAi[183]), .Y(
        b3_P_F_6_am_1));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[61]), .B(
        b11_OFWNT9L_8tZ[93]), .C(b4_nUAi[183]), .D(b4_nUAi[184]), .Y(
        b3_P_F_6_bm_1));
    
endmodule


module b8_1LbcQDr1_x_134_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [20:20] mdiclink_reg;
input  [134:134] b11_OFWNT9L_8tZ;
input  [62:60] b4_nUAi;
output [20:20] b6_2ZTGIf;

    wire b3_P_F_6_bm_85, b3_P_F_6_am_85, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_85), .B(
        b4_nUAi[62]), .C(b3_P_F_6_am_85), .Y(b6_2ZTGIf[20]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[20]), .B(
        b11_OFWNT9L_8tZ[134]), .C(b4_nUAi[61]), .D(b4_nUAi[60]), .Y(
        b3_P_F_6_am_85));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[20]), .B(
        b11_OFWNT9L_8tZ[134]), .C(b4_nUAi[60]), .D(b4_nUAi[61]), .Y(
        b3_P_F_6_bm_85));
    
endmodule


module b8_1LbcQDr1_x_94_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [60:60] mdiclink_reg;
input  [94:94] b11_OFWNT9L_8tZ;
input  [182:180] b4_nUAi;
output [60:60] b6_2ZTGIf;

    wire b3_P_F_6_bm_2, b3_P_F_6_am_2, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_2), .B(
        b4_nUAi[182]), .C(b3_P_F_6_am_2), .Y(b6_2ZTGIf[60]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[60]), .B(
        b11_OFWNT9L_8tZ[94]), .C(b4_nUAi[181]), .D(b4_nUAi[180]), .Y(
        b3_P_F_6_am_2));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[60]), .B(
        b11_OFWNT9L_8tZ[94]), .C(b4_nUAi[180]), .D(b4_nUAi[181]), .Y(
        b3_P_F_6_bm_2));
    
endmodule


module b8_1LbcQDr1_x_62_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [92:92] mdiclink_reg;
input  [62:62] b11_OFWNT9L_8tZ;
input  [278:276] b4_nUAi;
output [92:92] b6_2ZTGIf;

    wire b3_P_F_6_bm_22, b3_P_F_6_am_22, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_22), .B(
        b4_nUAi[278]), .C(b3_P_F_6_am_22), .Y(b6_2ZTGIf[92]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[92]), .B(
        b11_OFWNT9L_8tZ[62]), .C(b4_nUAi[277]), .D(b4_nUAi[276]), .Y(
        b3_P_F_6_am_22));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[92]), .B(
        b11_OFWNT9L_8tZ[62]), .C(b4_nUAi[276]), .D(b4_nUAi[277]), .Y(
        b3_P_F_6_bm_22));
    
endmodule


module b8_1LbcQDr1_x_78_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [76:76] mdiclink_reg;
input  [78:78] b11_OFWNT9L_8tZ;
input  [230:228] b4_nUAi;
output [76:76] b6_2ZTGIf;

    wire b3_P_F_6_bm_12, b3_P_F_6_am_12, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_12), .B(
        b4_nUAi[230]), .C(b3_P_F_6_am_12), .Y(b6_2ZTGIf[76]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[76]), .B(
        b11_OFWNT9L_8tZ[78]), .C(b4_nUAi[229]), .D(b4_nUAi[228]), .Y(
        b3_P_F_6_am_12));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[76]), .B(
        b11_OFWNT9L_8tZ[78]), .C(b4_nUAi[228]), .D(b4_nUAi[229]), .Y(
        b3_P_F_6_bm_12));
    
endmodule


module b8_1LbcQDr1_x_138_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [16:16] mdiclink_reg;
input  [138:138] b11_OFWNT9L_8tZ;
input  [49:48] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[16]), .B(
        b11_OFWNT9L_8tZ[138]), .C(b4_nUAi[49]), .D(b4_nUAi[48]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[16]), .B(
        b11_OFWNT9L_8tZ[138]), .C(b4_nUAi[49]), .D(b4_nUAi[48]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_117_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [37:37] mdiclink_reg;
input  [117:117] b11_OFWNT9L_8tZ;
input  [113:111] b4_nUAi;
output [37:37] b6_2ZTGIf;

    wire b3_P_F_6_bm_94, b3_P_F_6_am_94, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_94), .B(
        b4_nUAi[113]), .C(b3_P_F_6_am_94), .Y(b6_2ZTGIf[37]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[37]), .B(
        b11_OFWNT9L_8tZ[117]), .C(b4_nUAi[112]), .D(b4_nUAi[111]), .Y(
        b3_P_F_6_am_94));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[37]), .B(
        b11_OFWNT9L_8tZ[117]), .C(b4_nUAi[111]), .D(b4_nUAi[112]), .Y(
        b3_P_F_6_bm_94));
    
endmodule


module b8_1LbcQDr1_x_41_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [113:113] mdiclink_reg;
input  [41:41] b11_OFWNT9L_8tZ;
input  [340:339] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[113]), .B(
        b11_OFWNT9L_8tZ[41]), .C(b4_nUAi[340]), .D(b4_nUAi[339]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[113]), .B(
        b11_OFWNT9L_8tZ[41]), .C(b4_nUAi[340]), .D(b4_nUAi[339]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_66_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [88:88] mdiclink_reg;
input  [66:66] b11_OFWNT9L_8tZ;
input  [265:264] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[88]), .B(
        b11_OFWNT9L_8tZ[66]), .C(b4_nUAi[265]), .D(b4_nUAi[264]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[88]), .B(
        b11_OFWNT9L_8tZ[66]), .C(b4_nUAi[265]), .D(b4_nUAi[264]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_51_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [103:103] mdiclink_reg;
input  [51:51] b11_OFWNT9L_8tZ;
input  [311:309] b4_nUAi;
output [103:103] b6_2ZTGIf;

    wire b3_P_F_6_bm_35, b3_P_F_6_am_35, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_35), .B(
        b4_nUAi[311]), .C(b3_P_F_6_am_35), .Y(b6_2ZTGIf[103]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[103]), .B(
        b11_OFWNT9L_8tZ[51]), .C(b4_nUAi[310]), .D(b4_nUAi[309]), .Y(
        b3_P_F_6_am_35));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[103]), .B(
        b11_OFWNT9L_8tZ[51]), .C(b4_nUAi[309]), .D(b4_nUAi[310]), .Y(
        b3_P_F_6_bm_35));
    
endmodule


module b8_1LbcQDr1_x_98_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [56:56] mdiclink_reg;
input  [98:98] b11_OFWNT9L_8tZ;
input  [169:168] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[56]), .B(
        b11_OFWNT9L_8tZ[98]), .C(b4_nUAi[169]), .D(b4_nUAi[168]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[56]), .B(
        b11_OFWNT9L_8tZ[98]), .C(b4_nUAi[169]), .D(b4_nUAi[168]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_70_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [84:84] mdiclink_reg;
input  [70:70] b11_OFWNT9L_8tZ;
input  [254:252] b4_nUAi;
output [84:84] b6_2ZTGIf;

    wire b3_P_F_6_bm_28, b3_P_F_6_am_28, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_28), .B(
        b4_nUAi[254]), .C(b3_P_F_6_am_28), .Y(b6_2ZTGIf[84]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[84]), .B(
        b11_OFWNT9L_8tZ[70]), .C(b4_nUAi[253]), .D(b4_nUAi[252]), .Y(
        b3_P_F_6_am_28));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[84]), .B(
        b11_OFWNT9L_8tZ[70]), .C(b4_nUAi[252]), .D(b4_nUAi[253]), .Y(
        b3_P_F_6_bm_28));
    
endmodule


module b8_1LbcQDr1_x_2_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [152:152] mdiclink_reg;
input  [2:2] b11_OFWNT9L_8tZ;
input  [458:456] b4_nUAi;
output [152:152] b6_2ZTGIf;

    wire b3_P_F_6_bm_61, b3_P_F_6_am_61, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_61), .B(
        b4_nUAi[458]), .C(b3_P_F_6_am_61), .Y(b6_2ZTGIf[152]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[152]), .B(
        b11_OFWNT9L_8tZ[2]), .C(b4_nUAi[457]), .D(b4_nUAi[456]), .Y(
        b3_P_F_6_am_61));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[152]), .B(
        b11_OFWNT9L_8tZ[2]), .C(b4_nUAi[456]), .D(b4_nUAi[457]), .Y(
        b3_P_F_6_bm_61));
    
endmodule


module b8_1LbcQDr1_x_65_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [89:89] mdiclink_reg;
input  [65:65] b11_OFWNT9L_8tZ;
input  [269:267] b4_nUAi;
output [89:89] b6_2ZTGIf;

    wire b3_P_F_6_bm_24, b3_P_F_6_am_24, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_24), .B(
        b4_nUAi[269]), .C(b3_P_F_6_am_24), .Y(b6_2ZTGIf[89]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[89]), .B(
        b11_OFWNT9L_8tZ[65]), .C(b4_nUAi[268]), .D(b4_nUAi[267]), .Y(
        b3_P_F_6_am_24));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[89]), .B(
        b11_OFWNT9L_8tZ[65]), .C(b4_nUAi[267]), .D(b4_nUAi[268]), .Y(
        b3_P_F_6_bm_24));
    
endmodule


module b8_1LbcQDr1_x_153_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [1:1] mdiclink_reg;
input  [153:153] b11_OFWNT9L_8tZ;
input  [4:3] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[1]), .B(
        b11_OFWNT9L_8tZ[153]), .C(b4_nUAi[4]), .D(b4_nUAi[3]), .Y(N_27)
        );
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[1]), .B(
        b11_OFWNT9L_8tZ[153]), .C(b4_nUAi[4]), .D(b4_nUAi[3]), .Y(N_25)
        );
    
endmodule


module b8_1LbcQDr1_x_60_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [94:94] mdiclink_reg;
input  [60:60] b11_OFWNT9L_8tZ;
input  [284:282] b4_nUAi;
output [94:94] b6_2ZTGIf;

    wire b3_P_F_6_bm_20, b3_P_F_6_am_20, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_20), .B(
        b4_nUAi[284]), .C(b3_P_F_6_am_20), .Y(b6_2ZTGIf[94]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[94]), .B(
        b11_OFWNT9L_8tZ[60]), .C(b4_nUAi[283]), .D(b4_nUAi[282]), .Y(
        b3_P_F_6_am_20));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[94]), .B(
        b11_OFWNT9L_8tZ[60]), .C(b4_nUAi[282]), .D(b4_nUAi[283]), .Y(
        b3_P_F_6_bm_20));
    
endmodule


module b8_1LbcQDr1_x_32_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [122:122] mdiclink_reg;
input  [32:32] b11_OFWNT9L_8tZ;
input  [367:366] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[122]), .B(
        b11_OFWNT9L_8tZ[32]), .C(b4_nUAi[367]), .D(b4_nUAi[366]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[122]), .B(
        b11_OFWNT9L_8tZ[32]), .C(b4_nUAi[367]), .D(b4_nUAi[366]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_145_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [9:9] mdiclink_reg;
input  [145:145] b11_OFWNT9L_8tZ;
input  [29:27] b4_nUAi;
output [9:9] b6_2ZTGIf;

    wire b3_P_F_6_bm_71, b3_P_F_6_am_71, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_71), .B(
        b4_nUAi[29]), .C(b3_P_F_6_am_71), .Y(b6_2ZTGIf[9]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[9]), .B(
        b11_OFWNT9L_8tZ[145]), .C(b4_nUAi[28]), .D(b4_nUAi[27]), .Y(
        b3_P_F_6_am_71));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[9]), .B(
        b11_OFWNT9L_8tZ[145]), .C(b4_nUAi[27]), .D(b4_nUAi[28]), .Y(
        b3_P_F_6_bm_71));
    
endmodule


module b8_1LbcQDr1_x_126_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [28:28] mdiclink_reg;
input  [126:126] b11_OFWNT9L_8tZ;
input  [86:84] b4_nUAi;
output [28:28] b6_2ZTGIf;

    wire b3_P_F_6_bm_79, b3_P_F_6_am_79, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_79), .B(
        b4_nUAi[86]), .C(b3_P_F_6_am_79), .Y(b6_2ZTGIf[28]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[28]), .B(
        b11_OFWNT9L_8tZ[126]), .C(b4_nUAi[85]), .D(b4_nUAi[84]), .Y(
        b3_P_F_6_am_79));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[28]), .B(
        b11_OFWNT9L_8tZ[126]), .C(b4_nUAi[84]), .D(b4_nUAi[85]), .Y(
        b3_P_F_6_bm_79));
    
endmodule


module b8_1LbcQDr1_x_86_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [68:68] mdiclink_reg;
input  [86:86] b11_OFWNT9L_8tZ;
input  [206:204] b4_nUAi;
output [68:68] b6_2ZTGIf;

    wire b3_P_F_6_bm_18, b3_P_F_6_am_18, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_18), .B(
        b4_nUAi[206]), .C(b3_P_F_6_am_18), .Y(b6_2ZTGIf[68]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[68]), .B(
        b11_OFWNT9L_8tZ[86]), .C(b4_nUAi[205]), .D(b4_nUAi[204]), .Y(
        b3_P_F_6_am_18));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[68]), .B(
        b11_OFWNT9L_8tZ[86]), .C(b4_nUAi[204]), .D(b4_nUAi[205]), .Y(
        b3_P_F_6_bm_18));
    
endmodule


module b8_1LbcQDr1_x_57_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [97:97] mdiclink_reg;
input  [57:57] b11_OFWNT9L_8tZ;
input  [292:291] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[97]), .B(
        b11_OFWNT9L_8tZ[57]), .C(b4_nUAi[292]), .D(b4_nUAi[291]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[97]), .B(
        b11_OFWNT9L_8tZ[57]), .C(b4_nUAi[292]), .D(b4_nUAi[291]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_81_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [73:73] mdiclink_reg;
input  [81:81] b11_OFWNT9L_8tZ;
input  [221:219] b4_nUAi;
output [73:73] b6_2ZTGIf;

    wire b3_P_F_6_bm_14, b3_P_F_6_am_14, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_14), .B(
        b4_nUAi[221]), .C(b3_P_F_6_am_14), .Y(b6_2ZTGIf[73]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[73]), .B(
        b11_OFWNT9L_8tZ[81]), .C(b4_nUAi[220]), .D(b4_nUAi[219]), .Y(
        b3_P_F_6_am_14));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[73]), .B(
        b11_OFWNT9L_8tZ[81]), .C(b4_nUAi[219]), .D(b4_nUAi[220]), .Y(
        b3_P_F_6_bm_14));
    
endmodule


module b8_1LbcQDr1_x_141_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [13:13] mdiclink_reg;
input  [141:141] b11_OFWNT9L_8tZ;
input  [41:39] b4_nUAi;
output [13:13] b6_2ZTGIf;

    wire b3_P_F_6_bm_68, b3_P_F_6_am_68, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_68), .B(
        b4_nUAi[41]), .C(b3_P_F_6_am_68), .Y(b6_2ZTGIf[13]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[13]), .B(
        b11_OFWNT9L_8tZ[141]), .C(b4_nUAi[40]), .D(b4_nUAi[39]), .Y(
        b3_P_F_6_am_68));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[13]), .B(
        b11_OFWNT9L_8tZ[141]), .C(b4_nUAi[39]), .D(b4_nUAi[40]), .Y(
        b3_P_F_6_bm_68));
    
endmodule


module b8_1LbcQDr1_x_111_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [43:43] mdiclink_reg;
input  [111:111] b11_OFWNT9L_8tZ;
input  [131:129] b4_nUAi;
output [43:43] b6_2ZTGIf;

    wire b3_P_F_6_bm_90, b3_P_F_6_am_90, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_90), .B(
        b4_nUAi[131]), .C(b3_P_F_6_am_90), .Y(b6_2ZTGIf[43]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[43]), .B(
        b11_OFWNT9L_8tZ[111]), .C(b4_nUAi[130]), .D(b4_nUAi[129]), .Y(
        b3_P_F_6_am_90));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[43]), .B(
        b11_OFWNT9L_8tZ[111]), .C(b4_nUAi[129]), .D(b4_nUAi[130]), .Y(
        b3_P_F_6_bm_90));
    
endmodule


module b8_1LbcQDr1_x_29_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [125:125] mdiclink_reg;
input  [29:29] b11_OFWNT9L_8tZ;
input  [377:375] b4_nUAi;
output [125:125] b6_2ZTGIf;

    wire b3_P_F_6_bm_41, b3_P_F_6_am_41, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_41), .B(
        b4_nUAi[377]), .C(b3_P_F_6_am_41), .Y(b6_2ZTGIf[125]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[125]), .B(
        b11_OFWNT9L_8tZ[29]), .C(b4_nUAi[376]), .D(b4_nUAi[375]), .Y(
        b3_P_F_6_am_41));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[125]), .B(
        b11_OFWNT9L_8tZ[29]), .C(b4_nUAi[375]), .D(b4_nUAi[376]), .Y(
        b3_P_F_6_bm_41));
    
endmodule


module b8_1LbcQDr1_x_101_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [53:53] mdiclink_reg;
input  [101:101] b11_OFWNT9L_8tZ;
input  [161:159] b4_nUAi;
output [53:53] b6_2ZTGIf;

    wire b3_P_F_6_bm_7, b3_P_F_6_am_7, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_7), .B(
        b4_nUAi[161]), .C(b3_P_F_6_am_7), .Y(b6_2ZTGIf[53]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[53]), .B(
        b11_OFWNT9L_8tZ[101]), .C(b4_nUAi[160]), .D(b4_nUAi[159]), .Y(
        b3_P_F_6_am_7));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[53]), .B(
        b11_OFWNT9L_8tZ[101]), .C(b4_nUAi[159]), .D(b4_nUAi[160]), .Y(
        b3_P_F_6_bm_7));
    
endmodule


module b8_1LbcQDr1_x_125_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [29:29] mdiclink_reg;
input  [125:125] b11_OFWNT9L_8tZ;
input  [89:87] b4_nUAi;
output [29:29] b6_2ZTGIf;

    wire b3_P_F_6_bm_78, b3_P_F_6_am_78, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_78), .B(
        b4_nUAi[89]), .C(b3_P_F_6_am_78), .Y(b6_2ZTGIf[29]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[29]), .B(
        b11_OFWNT9L_8tZ[125]), .C(b4_nUAi[88]), .D(b4_nUAi[87]), .Y(
        b3_P_F_6_am_78));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[29]), .B(
        b11_OFWNT9L_8tZ[125]), .C(b4_nUAi[87]), .D(b4_nUAi[88]), .Y(
        b3_P_F_6_bm_78));
    
endmodule


module b8_1LbcQDr1_x_4_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [150:150] mdiclink_reg;
input  [4:4] b11_OFWNT9L_8tZ;
input  [451:450] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[150]), .B(
        b11_OFWNT9L_8tZ[4]), .C(b4_nUAi[451]), .D(b4_nUAi[450]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[150]), .B(
        b11_OFWNT9L_8tZ[4]), .C(b4_nUAi[451]), .D(b4_nUAi[450]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_85_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [69:69] mdiclink_reg;
input  [85:85] b11_OFWNT9L_8tZ;
input  [209:207] b4_nUAi;
output [69:69] b6_2ZTGIf;

    wire b3_P_F_6_bm_17, b3_P_F_6_am_17, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_17), .B(
        b4_nUAi[209]), .C(b3_P_F_6_am_17), .Y(b6_2ZTGIf[69]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[69]), .B(
        b11_OFWNT9L_8tZ[85]), .C(b4_nUAi[208]), .D(b4_nUAi[207]), .Y(
        b3_P_F_6_am_17));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[69]), .B(
        b11_OFWNT9L_8tZ[85]), .C(b4_nUAi[207]), .D(b4_nUAi[208]), .Y(
        b3_P_F_6_bm_17));
    
endmodule


module b8_1LbcQDr1_x_108_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [46:46] mdiclink_reg;
input  [108:108] b11_OFWNT9L_8tZ;
input  [140:138] b4_nUAi;
output [46:46] b6_2ZTGIf;

    wire b3_P_F_6_bm_87, b3_P_F_6_am_87, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_87), .B(
        b4_nUAi[140]), .C(b3_P_F_6_am_87), .Y(b6_2ZTGIf[46]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[46]), .B(
        b11_OFWNT9L_8tZ[108]), .C(b4_nUAi[139]), .D(b4_nUAi[138]), .Y(
        b3_P_F_6_am_87));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[46]), .B(
        b11_OFWNT9L_8tZ[108]), .C(b4_nUAi[138]), .D(b4_nUAi[139]), .Y(
        b3_P_F_6_bm_87));
    
endmodule


module b8_1LbcQDr1_x_25_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       N_27,
       N_25
    );
input  [129:129] mdiclink_reg;
input  [25:25] b11_OFWNT9L_8tZ;
input  [388:387] b4_nUAi;
output N_27;
output N_25;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8485) )  b3_P_F_5 (.A(mdiclink_reg[129]), .B(
        b11_OFWNT9L_8tZ[25]), .C(b4_nUAi[388]), .D(b4_nUAi[387]), .Y(
        N_27));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_3 (.A(mdiclink_reg[129]), .B(
        b11_OFWNT9L_8tZ[25]), .C(b4_nUAi[388]), .D(b4_nUAi[387]), .Y(
        N_25));
    
endmodule


module b8_1LbcQDr1_x_69_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b6_2ZTGIf
    );
input  [85:85] mdiclink_reg;
input  [69:69] b11_OFWNT9L_8tZ;
input  [257:255] b4_nUAi;
output [85:85] b6_2ZTGIf;

    wire b3_P_F_6_bm_27, b3_P_F_6_am_27, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hB8) )  b3_P_F_6_ns (.A(b3_P_F_6_bm_27), .B(
        b4_nUAi[257]), .C(b3_P_F_6_am_27), .Y(b6_2ZTGIf[85]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h12FA) )  b3_P_F_6_am (.A(mdiclink_reg[85]), .B(
        b11_OFWNT9L_8tZ[69]), .C(b4_nUAi[256]), .D(b4_nUAi[255]), .Y(
        b3_P_F_6_am_27));
    CFG4 #( .INIT(16'h8845) )  b3_P_F_6_bm (.A(mdiclink_reg[85]), .B(
        b11_OFWNT9L_8tZ[69]), .C(b4_nUAi[255]), .D(b4_nUAi[256]), .Y(
        b3_P_F_6_bm_27));
    
endmodule


module b11_PSyil9s1fkT_x(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b4_nUAi,
       b11_uUT0JC4gFrY,
       b7_PSyi3wy,
       BW_clk_c
    );
input  [154:0] mdiclink_reg;
input  [154:0] b11_OFWNT9L_8tZ;
input  [463:0] b4_nUAi;
output [1:1] b11_uUT0JC4gFrY;
input  b7_PSyi3wy;
input  BW_clk_c;

    wire N_27, N_25, N_27_0, N_25_0, N_27_1, N_25_1, N_27_2, N_25_2, 
        \b6_2ZTGIf[4] , \b6_2ZTGIf[5] , \b6_2ZTGIf[6] , \b6_2ZTGIf[7] , 
        N_27_3, N_25_3, \b6_2ZTGIf[9] , N_27_4, N_25_4, 
        \b6_2ZTGIf[11] , \b6_2ZTGIf[12] , \b6_2ZTGIf[13] , 
        \b6_2ZTGIf[14] , \b6_2ZTGIf[15] , N_27_5, N_25_5, N_27_6, 
        N_25_6, N_27_7, N_25_7, N_27_8, N_25_8, \b6_2ZTGIf[20] , 
        \b6_2ZTGIf[21] , \b6_2ZTGIf[22] , \b6_2ZTGIf[23] , N_27_9, 
        N_25_9, \b6_2ZTGIf[25] , N_27_10, N_25_10, \b6_2ZTGIf[27] , 
        \b6_2ZTGIf[28] , \b6_2ZTGIf[29] , \b6_2ZTGIf[30] , 
        \b6_2ZTGIf[31] , N_27_11, N_25_11, N_27_12, N_25_12, N_27_13, 
        N_25_13, N_27_14, N_25_14, \b6_2ZTGIf[36] , \b6_2ZTGIf[37] , 
        \b6_2ZTGIf[38] , \b6_2ZTGIf[39] , N_27_15, N_25_15, 
        \b6_2ZTGIf[41] , N_27_16, N_25_16, \b6_2ZTGIf[43] , 
        \b6_2ZTGIf[44] , \b6_2ZTGIf[45] , \b6_2ZTGIf[46] , 
        \b6_2ZTGIf[47] , N_27_17, N_25_17, N_27_18, N_25_18, N_27_19, 
        N_25_19, N_27_20, N_25_20, \b6_2ZTGIf[52] , \b6_2ZTGIf[53] , 
        \b6_2ZTGIf[54] , \b6_2ZTGIf[55] , N_27_21, N_25_21, 
        \b6_2ZTGIf[57] , N_27_22, N_25_22, \b6_2ZTGIf[59] , 
        \b6_2ZTGIf[60] , \b6_2ZTGIf[61] , \b6_2ZTGIf[62] , 
        \b6_2ZTGIf[63] , N_27_23, N_25_23, N_27_24, N_25_24, N_27_25, 
        N_25_25, N_27_26, N_25_26, \b6_2ZTGIf[68] , \b6_2ZTGIf[69] , 
        \b6_2ZTGIf[70] , \b6_2ZTGIf[71] , N_27_27, N_25_27, 
        \b6_2ZTGIf[73] , N_27_28, N_25_28, \b6_2ZTGIf[75] , 
        \b6_2ZTGIf[76] , \b6_2ZTGIf[77] , \b6_2ZTGIf[78] , 
        \b6_2ZTGIf[79] , N_27_29, N_25_29, N_27_30, N_25_30, N_27_31, 
        N_25_31, N_27_32, N_25_32, \b6_2ZTGIf[84] , \b6_2ZTGIf[85] , 
        \b6_2ZTGIf[86] , \b6_2ZTGIf[87] , N_27_33, N_25_33, 
        \b6_2ZTGIf[89] , N_27_34, N_25_34, \b6_2ZTGIf[91] , 
        \b6_2ZTGIf[92] , \b6_2ZTGIf[93] , \b6_2ZTGIf[94] , 
        \b6_2ZTGIf[95] , N_27_35, N_25_35, N_27_36, N_25_36, N_27_37, 
        N_25_37, N_27_38, N_25_38, \b6_2ZTGIf[100] , \b6_2ZTGIf[101] , 
        \b6_2ZTGIf[102] , \b6_2ZTGIf[103] , N_27_39, N_25_39, 
        \b6_2ZTGIf[105] , N_27_40, N_25_40, \b6_2ZTGIf[107] , 
        \b6_2ZTGIf[108] , \b6_2ZTGIf[109] , \b6_2ZTGIf[110] , 
        \b6_2ZTGIf[111] , N_27_41, N_25_41, N_27_42, N_25_42, N_27_43, 
        N_25_43, N_27_44, N_25_44, \b6_2ZTGIf[116] , \b6_2ZTGIf[117] , 
        \b6_2ZTGIf[118] , \b6_2ZTGIf[119] , N_27_45, N_25_45, 
        \b6_2ZTGIf[121] , N_27_46, N_25_46, \b6_2ZTGIf[123] , 
        \b6_2ZTGIf[124] , \b6_2ZTGIf[125] , \b6_2ZTGIf[126] , 
        \b6_2ZTGIf[127] , N_27_47, N_25_47, N_27_48, N_25_48, N_27_49, 
        N_25_49, N_27_50, N_25_50, \b6_2ZTGIf[132] , \b6_2ZTGIf[133] , 
        \b6_2ZTGIf[134] , \b6_2ZTGIf[135] , N_27_51, N_25_51, 
        \b6_2ZTGIf[137] , N_27_52, N_25_52, \b6_2ZTGIf[139] , 
        \b6_2ZTGIf[140] , \b6_2ZTGIf[141] , \b6_2ZTGIf[142] , 
        \b6_2ZTGIf[143] , \b6_2ZTGIf[144] , \b6_2ZTGIf[145] , N_27_53, 
        N_25_53, \b6_2ZTGIf[147] , N_27_54, N_25_54, \b6_2ZTGIf[149] , 
        N_27_55, N_25_55, N_27_56, N_25_56, \b6_2ZTGIf[152] , 
        \b6_2ZTGIf[153] , \b6_2ZTGIf[154] , GND_net_1, VCC_net_1;
    
    b8_1LbcQDr1_x_26_0 b9_1LbcgKGIS (.mdiclink_reg({mdiclink_reg[128]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[26]}), .b4_nUAi({
        b4_nUAi[385], b4_nUAi[384]}), .N_27(N_27_47), .N_25(N_25_47));
    b8_1LbcQDr1_x_80_0 b8_1LbcgKxQ0 (.mdiclink_reg({mdiclink_reg[74]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[80]}), .b4_nUAi({
        b4_nUAi[223], b4_nUAi[222]}), .N_27(N_27_28), .N_25(N_25_28));
    b8_1LbcQDr1_x_3_0 b9_1LbcgKGUn (.mdiclink_reg({mdiclink_reg[151]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[3]}), .b4_nUAi({b4_nUAi[454], 
        b4_nUAi[453]}), .N_27(N_27_56), .N_25(N_25_56));
    b8_1LbcQDr1_x_27_0 b9_1LbcgKGIe (.mdiclink_reg({mdiclink_reg[127]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[27]}), .b4_nUAi({
        b4_nUAi[383], b4_nUAi[382], b4_nUAi[381]}), .b6_2ZTGIf({
        \b6_2ZTGIf[127] }));
    b8_1LbcQDr1_x_140_0 b8_1LbcgKGQ0 (.mdiclink_reg({mdiclink_reg[14]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[140]}), .b4_nUAi({
        b4_nUAi[44], b4_nUAi[43], b4_nUAi[42]}), .b6_2ZTGIf({
        \b6_2ZTGIf[14] }));
    b8_1LbcQDr1_x_83_0 b8_1LbcgKxS (.mdiclink_reg({mdiclink_reg[71]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[83]}), .b4_nUAi({
        b4_nUAi[215], b4_nUAi[214], b4_nUAi[213]}), .b6_2ZTGIf({
        \b6_2ZTGIf[71] }));
    b8_1LbcQDr1_x_143_0 b8_1LbcgKGS (.mdiclink_reg({mdiclink_reg[11]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[143]}), .b4_nUAi({
        b4_nUAi[35], b4_nUAi[34], b4_nUAi[33]}), .b6_2ZTGIf({
        \b6_2ZTGIf[11] }));
    b8_1LbcQDr1_x_34_0 b9_1LbcgKGIm (.mdiclink_reg({mdiclink_reg[120]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[34]}), .b4_nUAi({
        b4_nUAi[361], b4_nUAi[360]}), .N_27(N_27_45), .N_25(N_25_45));
    b8_1LbcQDr1_x_84_0 b8_1LbcgKxR (.mdiclink_reg({mdiclink_reg[70]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[84]}), .b4_nUAi({
        b4_nUAi[212], b4_nUAi[211], b4_nUAi[210]}), .b6_2ZTGIf({
        \b6_2ZTGIf[70] }));
    b8_1LbcQDr1_x_144_0 b8_1LbcgKGR (.mdiclink_reg({mdiclink_reg[10]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[144]}), .b4_nUAi({
        b4_nUAi[31], b4_nUAi[30]}), .N_27(N_27_4), .N_25(N_25_4));
    b8_1LbcQDr1_x_103_0 b8_1LbcgKIS (.mdiclink_reg({mdiclink_reg[51]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[103]}), .b4_nUAi({
        b4_nUAi[154], b4_nUAi[153]}), .N_27(N_27_20), .N_25(N_25_20));
    b16_CRGcTCua_eH4_uui_x_0 b6_2ZGFQ9 (.b11_uUT0JC4gFrY({
        b11_uUT0JC4gFrY[1]}), .b6_2ZTGIf_3(\b6_2ZTGIf[7] ), 
        .b6_2ZTGIf_5(\b6_2ZTGIf[9] ), .b6_2ZTGIf_7(\b6_2ZTGIf[11] ), 
        .b6_2ZTGIf_8(\b6_2ZTGIf[12] ), .b6_2ZTGIf_9(\b6_2ZTGIf[13] ), 
        .b6_2ZTGIf_10(\b6_2ZTGIf[14] ), .b6_2ZTGIf_11(\b6_2ZTGIf[15] ), 
        .b6_2ZTGIf_2(\b6_2ZTGIf[6] ), .b6_2ZTGIf_1(\b6_2ZTGIf[5] ), 
        .b6_2ZTGIf_0(\b6_2ZTGIf[4] ), .b6_2ZTGIf_19(\b6_2ZTGIf[23] ), 
        .b6_2ZTGIf_21(\b6_2ZTGIf[25] ), .b6_2ZTGIf_23(\b6_2ZTGIf[27] ), 
        .b6_2ZTGIf_24(\b6_2ZTGIf[28] ), .b6_2ZTGIf_25(\b6_2ZTGIf[29] ), 
        .b6_2ZTGIf_26(\b6_2ZTGIf[30] ), .b6_2ZTGIf_27(\b6_2ZTGIf[31] ), 
        .b6_2ZTGIf_18(\b6_2ZTGIf[22] ), .b6_2ZTGIf_17(\b6_2ZTGIf[21] ), 
        .b6_2ZTGIf_16(\b6_2ZTGIf[20] ), .b6_2ZTGIf_35(\b6_2ZTGIf[39] ), 
        .b6_2ZTGIf_37(\b6_2ZTGIf[41] ), .b6_2ZTGIf_39(\b6_2ZTGIf[43] ), 
        .b6_2ZTGIf_40(\b6_2ZTGIf[44] ), .b6_2ZTGIf_41(\b6_2ZTGIf[45] ), 
        .b6_2ZTGIf_42(\b6_2ZTGIf[46] ), .b6_2ZTGIf_43(\b6_2ZTGIf[47] ), 
        .b6_2ZTGIf_34(\b6_2ZTGIf[38] ), .b6_2ZTGIf_33(\b6_2ZTGIf[37] ), 
        .b6_2ZTGIf_32(\b6_2ZTGIf[36] ), .b6_2ZTGIf_51(\b6_2ZTGIf[55] ), 
        .b6_2ZTGIf_53(\b6_2ZTGIf[57] ), .b6_2ZTGIf_55(\b6_2ZTGIf[59] ), 
        .b6_2ZTGIf_56(\b6_2ZTGIf[60] ), .b6_2ZTGIf_57(\b6_2ZTGIf[61] ), 
        .b6_2ZTGIf_58(\b6_2ZTGIf[62] ), .b6_2ZTGIf_59(\b6_2ZTGIf[63] ), 
        .b6_2ZTGIf_50(\b6_2ZTGIf[54] ), .b6_2ZTGIf_49(\b6_2ZTGIf[53] ), 
        .b6_2ZTGIf_48(\b6_2ZTGIf[52] ), .b6_2ZTGIf_67(\b6_2ZTGIf[71] ), 
        .b6_2ZTGIf_69(\b6_2ZTGIf[73] ), .b6_2ZTGIf_71(\b6_2ZTGIf[75] ), 
        .b6_2ZTGIf_72(\b6_2ZTGIf[76] ), .b6_2ZTGIf_73(\b6_2ZTGIf[77] ), 
        .b6_2ZTGIf_74(\b6_2ZTGIf[78] ), .b6_2ZTGIf_75(\b6_2ZTGIf[79] ), 
        .b6_2ZTGIf_66(\b6_2ZTGIf[70] ), .b6_2ZTGIf_65(\b6_2ZTGIf[69] ), 
        .b6_2ZTGIf_64(\b6_2ZTGIf[68] ), .b6_2ZTGIf_83(\b6_2ZTGIf[87] ), 
        .b6_2ZTGIf_85(\b6_2ZTGIf[89] ), .b6_2ZTGIf_87(\b6_2ZTGIf[91] ), 
        .b6_2ZTGIf_88(\b6_2ZTGIf[92] ), .b6_2ZTGIf_89(\b6_2ZTGIf[93] ), 
        .b6_2ZTGIf_90(\b6_2ZTGIf[94] ), .b6_2ZTGIf_91(\b6_2ZTGIf[95] ), 
        .b6_2ZTGIf_82(\b6_2ZTGIf[86] ), .b6_2ZTGIf_81(\b6_2ZTGIf[85] ), 
        .b6_2ZTGIf_80(\b6_2ZTGIf[84] ), .b6_2ZTGIf_99(\b6_2ZTGIf[103] )
        , .b6_2ZTGIf_101(\b6_2ZTGIf[105] ), .b6_2ZTGIf_103(
        \b6_2ZTGIf[107] ), .b6_2ZTGIf_104(\b6_2ZTGIf[108] ), 
        .b6_2ZTGIf_105(\b6_2ZTGIf[109] ), .b6_2ZTGIf_106(
        \b6_2ZTGIf[110] ), .b6_2ZTGIf_107(\b6_2ZTGIf[111] ), 
        .b6_2ZTGIf_98(\b6_2ZTGIf[102] ), .b6_2ZTGIf_97(
        \b6_2ZTGIf[101] ), .b6_2ZTGIf_96(\b6_2ZTGIf[100] ), 
        .b6_2ZTGIf_115(\b6_2ZTGIf[119] ), .b6_2ZTGIf_117(
        \b6_2ZTGIf[121] ), .b6_2ZTGIf_119(\b6_2ZTGIf[123] ), 
        .b6_2ZTGIf_120(\b6_2ZTGIf[124] ), .b6_2ZTGIf_121(
        \b6_2ZTGIf[125] ), .b6_2ZTGIf_122(\b6_2ZTGIf[126] ), 
        .b6_2ZTGIf_123(\b6_2ZTGIf[127] ), .b6_2ZTGIf_114(
        \b6_2ZTGIf[118] ), .b6_2ZTGIf_113(\b6_2ZTGIf[117] ), 
        .b6_2ZTGIf_112(\b6_2ZTGIf[116] ), .b6_2ZTGIf_131(
        \b6_2ZTGIf[135] ), .b6_2ZTGIf_133(\b6_2ZTGIf[137] ), 
        .b6_2ZTGIf_135(\b6_2ZTGIf[139] ), .b6_2ZTGIf_136(
        \b6_2ZTGIf[140] ), .b6_2ZTGIf_137(\b6_2ZTGIf[141] ), 
        .b6_2ZTGIf_138(\b6_2ZTGIf[142] ), .b6_2ZTGIf_139(
        \b6_2ZTGIf[143] ), .b6_2ZTGIf_130(\b6_2ZTGIf[134] ), 
        .b6_2ZTGIf_129(\b6_2ZTGIf[133] ), .b6_2ZTGIf_128(
        \b6_2ZTGIf[132] ), .b6_2ZTGIf_141(\b6_2ZTGIf[145] ), 
        .b6_2ZTGIf_143(\b6_2ZTGIf[147] ), .b6_2ZTGIf_145(
        \b6_2ZTGIf[149] ), .b6_2ZTGIf_150(\b6_2ZTGIf[154] ), 
        .b6_2ZTGIf_149(\b6_2ZTGIf[153] ), .b6_2ZTGIf_148(
        \b6_2ZTGIf[152] ), .b6_2ZTGIf_140(\b6_2ZTGIf[144] ), 
        .b4_nUAi_24(b4_nUAi[26]), .b4_nUAi_30(b4_nUAi[32]), .b4_nUAi_0(
        b4_nUAi[2]), .b4_nUAi_3(b4_nUAi[5]), .b4_nUAi_6(b4_nUAi[8]), 
        .b4_nUAi_9(b4_nUAi[11]), .b4_nUAi_72(b4_nUAi[74]), .b4_nUAi_78(
        b4_nUAi[80]), .b4_nUAi_48(b4_nUAi[50]), .b4_nUAi_51(
        b4_nUAi[53]), .b4_nUAi_54(b4_nUAi[56]), .b4_nUAi_57(
        b4_nUAi[59]), .b4_nUAi_120(b4_nUAi[122]), .b4_nUAi_126(
        b4_nUAi[128]), .b4_nUAi_96(b4_nUAi[98]), .b4_nUAi_99(
        b4_nUAi[101]), .b4_nUAi_102(b4_nUAi[104]), .b4_nUAi_105(
        b4_nUAi[107]), .b4_nUAi_168(b4_nUAi[170]), .b4_nUAi_174(
        b4_nUAi[176]), .b4_nUAi_144(b4_nUAi[146]), .b4_nUAi_147(
        b4_nUAi[149]), .b4_nUAi_150(b4_nUAi[152]), .b4_nUAi_153(
        b4_nUAi[155]), .b4_nUAi_216(b4_nUAi[218]), .b4_nUAi_222(
        b4_nUAi[224]), .b4_nUAi_192(b4_nUAi[194]), .b4_nUAi_195(
        b4_nUAi[197]), .b4_nUAi_198(b4_nUAi[200]), .b4_nUAi_201(
        b4_nUAi[203]), .b4_nUAi_264(b4_nUAi[266]), .b4_nUAi_270(
        b4_nUAi[272]), .b4_nUAi_240(b4_nUAi[242]), .b4_nUAi_243(
        b4_nUAi[245]), .b4_nUAi_246(b4_nUAi[248]), .b4_nUAi_249(
        b4_nUAi[251]), .b4_nUAi_312(b4_nUAi[314]), .b4_nUAi_318(
        b4_nUAi[320]), .b4_nUAi_288(b4_nUAi[290]), .b4_nUAi_291(
        b4_nUAi[293]), .b4_nUAi_294(b4_nUAi[296]), .b4_nUAi_297(
        b4_nUAi[299]), .b4_nUAi_360(b4_nUAi[362]), .b4_nUAi_366(
        b4_nUAi[368]), .b4_nUAi_336(b4_nUAi[338]), .b4_nUAi_339(
        b4_nUAi[341]), .b4_nUAi_342(b4_nUAi[344]), .b4_nUAi_345(
        b4_nUAi[347]), .b4_nUAi_408(b4_nUAi[410]), .b4_nUAi_414(
        b4_nUAi[416]), .b4_nUAi_384(b4_nUAi[386]), .b4_nUAi_387(
        b4_nUAi[389]), .b4_nUAi_390(b4_nUAi[392]), .b4_nUAi_393(
        b4_nUAi[395]), .b4_nUAi_438(b4_nUAi[440]), .b4_nUAi_444(
        b4_nUAi[446]), .b4_nUAi_450(b4_nUAi[452]), .b4_nUAi_453(
        b4_nUAi[455]), .BW_clk_c(BW_clk_c), .N_25(N_25_3), .N_27(
        N_27_3), .N_25_0(N_25_4), .N_27_0(N_27_4), .N_25_1(N_25), 
        .N_27_1(N_27), .N_25_2(N_25_0), .N_27_2(N_27_0), .N_25_3(
        N_25_1), .N_27_3(N_27_1), .N_25_4(N_25_2), .N_27_4(N_27_2), 
        .N_25_5(N_25_9), .N_27_5(N_27_9), .N_25_6(N_25_10), .N_27_6(
        N_27_10), .N_25_7(N_25_5), .N_27_7(N_27_5), .N_25_8(N_25_6), 
        .N_27_8(N_27_6), .N_25_9(N_25_7), .N_27_9(N_27_7), .N_25_10(
        N_25_8), .N_27_10(N_27_8), .N_25_11(N_25_15), .N_27_11(N_27_15)
        , .N_25_12(N_25_16), .N_27_12(N_27_16), .N_25_13(N_25_11), 
        .N_27_13(N_27_11), .N_25_14(N_25_12), .N_27_14(N_27_12), 
        .N_25_15(N_25_13), .N_27_15(N_27_13), .N_25_16(N_25_14), 
        .N_27_16(N_27_14), .N_25_17(N_25_21), .N_27_17(N_27_21), 
        .N_25_18(N_25_22), .N_27_18(N_27_22), .N_25_19(N_25_17), 
        .N_27_19(N_27_17), .N_25_20(N_25_18), .N_27_20(N_27_18), 
        .N_25_21(N_25_19), .N_27_21(N_27_19), .N_25_22(N_25_20), 
        .N_27_22(N_27_20), .N_25_23(N_25_27), .N_27_23(N_27_27), 
        .N_25_24(N_25_28), .N_27_24(N_27_28), .N_25_25(N_25_23), 
        .N_27_25(N_27_23), .N_25_26(N_25_24), .N_27_26(N_27_24), 
        .N_25_27(N_25_25), .N_27_27(N_27_25), .N_25_28(N_25_26), 
        .N_27_28(N_27_26), .N_25_29(N_25_33), .N_27_29(N_27_33), 
        .N_25_30(N_25_34), .N_27_30(N_27_34), .N_25_31(N_25_29), 
        .N_27_31(N_27_29), .N_25_32(N_25_30), .N_27_32(N_27_30), 
        .N_25_33(N_25_31), .N_27_33(N_27_31), .N_25_34(N_25_32), 
        .N_27_34(N_27_32), .N_25_35(N_25_39), .N_27_35(N_27_39), 
        .N_25_36(N_25_40), .N_27_36(N_27_40), .N_25_37(N_25_35), 
        .N_27_37(N_27_35), .N_25_38(N_25_36), .N_27_38(N_27_36), 
        .N_25_39(N_25_37), .N_27_39(N_27_37), .N_25_40(N_25_38), 
        .N_27_40(N_27_38), .N_25_41(N_25_45), .N_27_41(N_27_45), 
        .N_25_42(N_25_46), .N_27_42(N_27_46), .N_25_43(N_25_41), 
        .N_27_43(N_27_41), .N_25_44(N_25_42), .N_27_44(N_27_42), 
        .N_25_45(N_25_43), .N_27_45(N_27_43), .N_25_46(N_25_44), 
        .N_27_46(N_27_44), .N_25_47(N_25_51), .N_27_47(N_27_51), 
        .N_25_48(N_25_52), .N_27_48(N_27_52), .N_25_49(N_25_47), 
        .N_27_49(N_27_47), .N_25_50(N_25_48), .N_27_50(N_27_48), 
        .N_25_51(N_25_49), .N_27_51(N_27_49), .N_25_52(N_25_50), 
        .N_27_52(N_27_50), .N_25_53(N_25_53), .N_27_53(N_27_53), 
        .N_25_54(N_25_54), .N_27_54(N_27_54), .N_25_55(N_25_55), 
        .N_27_55(N_27_55), .N_25_56(N_25_56), .N_27_56(N_27_56));
    b8_1LbcQDr1_x_104_0 b8_1LbcgKIR (.mdiclink_reg({mdiclink_reg[50]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[104]}), .b4_nUAi({
        b4_nUAi[151], b4_nUAi[150]}), .N_27(N_27_19), .N_25(N_25_19));
    b8_1LbcQDr1_x_72_0 b8_1LbcgKbI (.mdiclink_reg({mdiclink_reg[82]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[72]}), .b4_nUAi({
        b4_nUAi[247], b4_nUAi[246]}), .N_27(N_27_31), .N_25(N_25_31));
    b8_1LbcQDr1_x_33_0 b9_1LbcgKGIn (.mdiclink_reg({mdiclink_reg[121]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[33]}), .b4_nUAi({
        b4_nUAi[365], b4_nUAi[364], b4_nUAi[363]}), .b6_2ZTGIf({
        \b6_2ZTGIf[121] }));
    b8_1LbcQDr1_x_129_0 b8_1LbcgKwU (.mdiclink_reg({mdiclink_reg[25]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[129]}), .b4_nUAi({
        b4_nUAi[77], b4_nUAi[76], b4_nUAi[75]}), .b6_2ZTGIf({
        \b6_2ZTGIf[25] }));
    b8_1LbcQDr1_x_89_0 b8_1LbcgKoU (.mdiclink_reg({mdiclink_reg[65]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[89]}), .b4_nUAi({
        b4_nUAi[196], b4_nUAi[195]}), .N_27(N_27_24), .N_25(N_25_24));
    b8_1LbcQDr1_x_120_0 b8_1LbcgKeQ0 (.mdiclink_reg({mdiclink_reg[34]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[120]}), .b4_nUAi({
        b4_nUAi[103], b4_nUAi[102]}), .N_27(N_27_13), .N_25(N_25_13));
    b8_1LbcQDr1_x_90_0 b8_1LbcgKoQ0 (.mdiclink_reg({mdiclink_reg[64]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[90]}), .b4_nUAi({
        b4_nUAi[193], b4_nUAi[192]}), .N_27(N_27_23), .N_25(N_25_23));
    b8_1LbcQDr1_x_10_0 b9_1LbcgKGQl0 (.mdiclink_reg({mdiclink_reg[144]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[10]}), .b4_nUAi({
        b4_nUAi[434], b4_nUAi[433], b4_nUAi[432]}), .b6_2ZTGIf({
        \b6_2ZTGIf[144] }));
    b8_1LbcQDr1_x_8_0 b9_1LbcgKGQ50 (.mdiclink_reg({mdiclink_reg[146]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[8]}), .b4_nUAi({
        b4_nUAi[439], b4_nUAi[438]}), .N_27(N_27_53), .N_25(N_25_53));
    b8_1LbcQDr1_x_1_0 b9_1LbcgKGUV (.mdiclink_reg({mdiclink_reg[153]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[1]}), .b4_nUAi({b4_nUAi[461], 
        b4_nUAi[460], b4_nUAi[459]}), .b6_2ZTGIf({\b6_2ZTGIf[153] }));
    b8_1LbcQDr1_x_130_0 b8_1LbcgKwQ0 (.mdiclink_reg({mdiclink_reg[24]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[130]}), .b4_nUAi({
        b4_nUAi[73], b4_nUAi[72]}), .N_27(N_27_9), .N_25(N_25_9));
    b8_1LbcQDr1_x_132_0 b8_1LbcgKwI (.mdiclink_reg({mdiclink_reg[22]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[132]}), .b4_nUAi({
        b4_nUAi[68], b4_nUAi[67], b4_nUAi[66]}), .b6_2ZTGIf({
        \b6_2ZTGIf[22] }));
    b8_1LbcQDr1_x_92_0 b8_1LbcgKoI (.mdiclink_reg({mdiclink_reg[62]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[92]}), .b4_nUAi({
        b4_nUAi[188], b4_nUAi[187], b4_nUAi[186]}), .b6_2ZTGIf({
        \b6_2ZTGIf[62] }));
    b8_1LbcQDr1_x_113_0 b8_1LbcgKES0 (.mdiclink_reg({mdiclink_reg[41]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[113]}), .b4_nUAi({
        b4_nUAi[125], b4_nUAi[124], b4_nUAi[123]}), .b6_2ZTGIf({
        \b6_2ZTGIf[41] }));
    b8_1LbcQDr1_x_76_0 b8_1LbcgKxn (.mdiclink_reg({mdiclink_reg[78]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[76]}), .b4_nUAi({
        b4_nUAi[236], b4_nUAi[235], b4_nUAi[234]}), .b6_2ZTGIf({
        \b6_2ZTGIf[78] }));
    b8_1LbcQDr1_x_136_0 b8_1LbcgKGn (.mdiclink_reg({mdiclink_reg[18]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[136]}), .b4_nUAi({
        b4_nUAi[55], b4_nUAi[54]}), .N_27(N_27_7), .N_25(N_25_7));
    b8_1LbcQDr1_x_67_0 b8_1LbcgKbJ (.mdiclink_reg({mdiclink_reg[87]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[67]}), .b4_nUAi({
        b4_nUAi[263], b4_nUAi[262], b4_nUAi[261]}), .b6_2ZTGIf({
        \b6_2ZTGIf[87] }));
    b8_1LbcQDr1_x_114_0 b8_1LbcgKER0 (.mdiclink_reg({mdiclink_reg[40]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[114]}), .b4_nUAi({
        b4_nUAi[121], b4_nUAi[120]}), .N_27(N_27_15), .N_25(N_25_15));
    b8_1LbcQDr1_x_118_0 b8_1LbcgKeA (.mdiclink_reg({mdiclink_reg[36]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[118]}), .b4_nUAi({
        b4_nUAi[110], b4_nUAi[109], b4_nUAi[108]}), .b6_2ZTGIf({
        \b6_2ZTGIf[36] }));
    b8_1LbcQDr1_x_96_0 b8_1LbcgKIn (.mdiclink_reg({mdiclink_reg[58]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[96]}), .b4_nUAi({
        b4_nUAi[175], b4_nUAi[174]}), .N_27(N_27_22), .N_25(N_25_22));
    b8_1LbcQDr1_x_31_0 b9_1LbcgKGIV (.mdiclink_reg({mdiclink_reg[123]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[31]}), .b4_nUAi({
        b4_nUAi[371], b4_nUAi[370], b4_nUAi[369]}), .b6_2ZTGIf({
        \b6_2ZTGIf[123] }));
    GND GND (.Y(GND_net_1));
    b8_1LbcQDr1_x_75_0 b8_1LbcgKxV (.mdiclink_reg({mdiclink_reg[79]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[75]}), .b4_nUAi({
        b4_nUAi[239], b4_nUAi[238], b4_nUAi[237]}), .b6_2ZTGIf({
        \b6_2ZTGIf[79] }));
    b8_1LbcQDr1_x_135_0 b8_1LbcgKGV (.mdiclink_reg({mdiclink_reg[19]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[135]}), .b4_nUAi({
        b4_nUAi[58], b4_nUAi[57]}), .N_27(N_27_8), .N_25(N_25_8));
    b8_1LbcQDr1_x_20_0 b9_1LbcgKGql (.mdiclink_reg({mdiclink_reg[134]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[20]}), .b4_nUAi({
        b4_nUAi[404], b4_nUAi[403], b4_nUAi[402]}), .b6_2ZTGIf({
        \b6_2ZTGIf[134] }));
    b8_1LbcQDr1_x_95_0 b8_1LbcgKIV (.mdiclink_reg({mdiclink_reg[59]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[95]}), .b4_nUAi({
        b4_nUAi[179], b4_nUAi[178], b4_nUAi[177]}), .b6_2ZTGIf({
        \b6_2ZTGIf[59] }));
    b8_1LbcQDr1_x_150_0 b7_1LbcgKE0 (.mdiclink_reg({mdiclink_reg[4]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[150]}), .b4_nUAi({
        b4_nUAi[14], b4_nUAi[13], b4_nUAi[12]}), .b6_2ZTGIf({
        \b6_2ZTGIf[4] }));
    b8_1LbcQDr1_x_18_0 b9_1LbcgKGq5 (.mdiclink_reg({mdiclink_reg[136]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[18]}), .b4_nUAi({
        b4_nUAi[409], b4_nUAi[408]}), .N_27(N_27_51), .N_25(N_25_51));
    b8_1LbcQDr1_x_127_0 b8_1LbcgKwJ (.mdiclink_reg({mdiclink_reg[27]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[127]}), .b4_nUAi({
        b4_nUAi[83], b4_nUAi[82], b4_nUAi[81]}), .b6_2ZTGIf({
        \b6_2ZTGIf[27] }));
    b8_1LbcQDr1_x_87_0 b8_1LbcgKoJ (.mdiclink_reg({mdiclink_reg[67]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[87]}), .b4_nUAi({
        b4_nUAi[202], b4_nUAi[201]}), .N_27(N_27_26), .N_25(N_25_26));
    b8_1LbcQDr1_x_40_0 b9_1LbcgKGSl (.mdiclink_reg({mdiclink_reg[114]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[40]}), .b4_nUAi({
        b4_nUAi[343], b4_nUAi[342]}), .N_27(N_27_43), .N_25(N_25_43));
    b8_1LbcQDr1_x_58_0 b8_1LbcgKJA (.mdiclink_reg({mdiclink_reg[96]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[58]}), .b4_nUAi({
        b4_nUAi[289], b4_nUAi[288]}), .N_27(N_27_35), .N_25(N_25_35));
    b8_1LbcQDr1_x_38_0 b9_1LbcgKGS5 (.mdiclink_reg({mdiclink_reg[116]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[38]}), .b4_nUAi({
        b4_nUAi[350], b4_nUAi[349], b4_nUAi[348]}), .b6_2ZTGIf({
        \b6_2ZTGIf[116] }));
    b8_1LbcQDr1_x_50_0 b9_1LbcgKGRl (.mdiclink_reg({mdiclink_reg[104]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[50]}), .b4_nUAi({
        b4_nUAi[313], b4_nUAi[312]}), .N_27(N_27_39), .N_25(N_25_39));
    b8_1LbcQDr1_x_121_0 b8_1LbcgKeq (.mdiclink_reg({mdiclink_reg[33]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[121]}), .b4_nUAi({
        b4_nUAi[100], b4_nUAi[99]}), .N_27(N_27_12), .N_25(N_25_12));
    b8_1LbcQDr1_x_48_0 b9_1LbcgKGR5 (.mdiclink_reg({mdiclink_reg[106]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[48]}), .b4_nUAi({
        b4_nUAi[319], b4_nUAi[318]}), .N_27(N_27_40), .N_25(N_25_40));
    b8_1LbcQDr1_x_106_0 b8_1LbcgKEn0 (.mdiclink_reg({mdiclink_reg[48]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[106]}), .b4_nUAi({
        b4_nUAi[145], b4_nUAi[144]}), .N_27(N_27_17), .N_25(N_25_17));
    b8_1LbcQDr1_x_79_0 b8_1LbcgKxU (.mdiclink_reg({mdiclink_reg[75]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[79]}), .b4_nUAi({
        b4_nUAi[227], b4_nUAi[226], b4_nUAi[225]}), .b6_2ZTGIf({
        \b6_2ZTGIf[75] }));
    b8_1LbcQDr1_x_139_0 b8_1LbcgKGU (.mdiclink_reg({mdiclink_reg[15]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[139]}), .b4_nUAi({
        b4_nUAi[47], b4_nUAi[46], b4_nUAi[45]}), .b6_2ZTGIf({
        \b6_2ZTGIf[15] }));
    b8_1LbcQDr1_x_147_0 b7_1LbcgKx (.mdiclink_reg({mdiclink_reg[7]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[147]}), .b4_nUAi({
        b4_nUAi[23], b4_nUAi[22], b4_nUAi[21]}), .b6_2ZTGIf({
        \b6_2ZTGIf[7] }));
    b8_1LbcQDr1_x_99_0 b8_1LbcgKIU (.mdiclink_reg({mdiclink_reg[55]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[99]}), .b4_nUAi({
        b4_nUAi[167], b4_nUAi[166], b4_nUAi[165]}), .b6_2ZTGIf({
        \b6_2ZTGIf[55] }));
    b8_1LbcQDr1_x_105_0 b8_1LbcgKEV0 (.mdiclink_reg({mdiclink_reg[49]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[105]}), .b4_nUAi({
        b4_nUAi[148], b4_nUAi[147]}), .N_27(N_27_18), .N_25(N_25_18));
    VCC VCC (.Y(VCC_net_1));
    b8_1LbcQDr1_x_110_0 b8_1LbcgKEQ0 (.mdiclink_reg({mdiclink_reg[44]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[110]}), .b4_nUAi({
        b4_nUAi[134], b4_nUAi[133], b4_nUAi[132]}), .b6_2ZTGIf({
        \b6_2ZTGIf[44] }));
    b8_1LbcQDr1_x_123_0 b8_1LbcgKeS (.mdiclink_reg({mdiclink_reg[31]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[123]}), .b4_nUAi({
        b4_nUAi[95], b4_nUAi[94], b4_nUAi[93]}), .b6_2ZTGIf({
        \b6_2ZTGIf[31] }));
    b8_1LbcQDr1_x_82_0 b8_1LbcgKxI (.mdiclink_reg({mdiclink_reg[72]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[82]}), .b4_nUAi({
        b4_nUAi[217], b4_nUAi[216]}), .N_27(N_27_27), .N_25(N_25_27));
    b8_1LbcQDr1_x_142_0 b8_1LbcgKGI (.mdiclink_reg({mdiclink_reg[12]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[142]}), .b4_nUAi({
        b4_nUAi[38], b4_nUAi[37], b4_nUAi[36]}), .b6_2ZTGIf({
        \b6_2ZTGIf[12] }));
    b8_1LbcQDr1_x_124_0 b8_1LbcgKeR (.mdiclink_reg({mdiclink_reg[30]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[124]}), .b4_nUAi({
        b4_nUAi[92], b4_nUAi[91], b4_nUAi[90]}), .b6_2ZTGIf({
        \b6_2ZTGIf[30] }));
    b8_1LbcQDr1_x_102_0 b8_1LbcgKII (.mdiclink_reg({mdiclink_reg[52]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[102]}), .b4_nUAi({
        b4_nUAi[158], b4_nUAi[157], b4_nUAi[156]}), .b6_2ZTGIf({
        \b6_2ZTGIf[52] }));
    b8_1LbcQDr1_x_12_0 b9_1LbcgKGQd0 (.mdiclink_reg({mdiclink_reg[142]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[12]}), .b4_nUAi({
        b4_nUAi[428], b4_nUAi[427], b4_nUAi[426]}), .b6_2ZTGIf({
        \b6_2ZTGIf[142] }));
    b8_1LbcQDr1_x_61_0 b8_1LbcgKJq (.mdiclink_reg({mdiclink_reg[93]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[61]}), .b4_nUAi({
        b4_nUAi[281], b4_nUAi[280], b4_nUAi[279]}), .b6_2ZTGIf({
        \b6_2ZTGIf[93] }));
    b8_1LbcQDr1_x_148_0 b7_1LbcgKo (.mdiclink_reg({mdiclink_reg[6]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[148]}), .b4_nUAi({
        b4_nUAi[20], b4_nUAi[19], b4_nUAi[18]}), .b6_2ZTGIf({
        \b6_2ZTGIf[6] }));
    b8_1LbcQDr1_x_9_0 b9_1LbcgKGQp0 (.mdiclink_reg({mdiclink_reg[145]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[9]}), .b4_nUAi({
        b4_nUAi[437], b4_nUAi[436], b4_nUAi[435]}), .b6_2ZTGIf({
        \b6_2ZTGIf[145] }));
    b8_1LbcQDr1_x_109_0 b8_1LbcgKEU0 (.mdiclink_reg({mdiclink_reg[45]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[109]}), .b4_nUAi({
        b4_nUAi[137], b4_nUAi[136], b4_nUAi[135]}), .b6_2ZTGIf({
        \b6_2ZTGIf[45] }));
    b8_1LbcQDr1_x_5_0 b9_1LbcgKGQq0 (.mdiclink_reg({mdiclink_reg[149]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[5]}), .b4_nUAi({
        b4_nUAi[449], b4_nUAi[448], b4_nUAi[447]}), .b6_2ZTGIf({
        \b6_2ZTGIf[149] }));
    b8_1LbcQDr1_x_63_0 b8_1LbcgKJS (.mdiclink_reg({mdiclink_reg[91]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[63]}), .b4_nUAi({
        b4_nUAi[275], b4_nUAi[274], b4_nUAi[273]}), .b6_2ZTGIf({
        \b6_2ZTGIf[91] }));
    b8_1LbcQDr1_x_149_0 b7_1LbcgKI (.mdiclink_reg({mdiclink_reg[5]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[149]}), .b4_nUAi({
        b4_nUAi[17], b4_nUAi[16], b4_nUAi[15]}), .b6_2ZTGIf({
        \b6_2ZTGIf[5] }));
    b8_1LbcQDr1_x_6_0 b9_1LbcgKGQS0 (.mdiclink_reg({mdiclink_reg[148]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[6]}), .b4_nUAi({
        b4_nUAi[445], b4_nUAi[444]}), .N_27(N_27_54), .N_25(N_25_54));
    b8_1LbcQDr1_x_64_0 b8_1LbcgKJR (.mdiclink_reg({mdiclink_reg[90]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[64]}), .b4_nUAi({
        b4_nUAi[271], b4_nUAi[270]}), .N_27(N_27_34), .N_25(N_25_34));
    b8_1LbcQDr1_x_22_0 b9_1LbcgKGqd (.mdiclink_reg({mdiclink_reg[132]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[22]}), .b4_nUAi({
        b4_nUAi[398], b4_nUAi[397], b4_nUAi[396]}), .b6_2ZTGIf({
        \b6_2ZTGIf[132] }));
    b8_1LbcQDr1_x_7_0 b9_1LbcgKGQe0 (.mdiclink_reg({mdiclink_reg[147]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[7]}), .b4_nUAi({
        b4_nUAi[443], b4_nUAi[442], b4_nUAi[441]}), .b6_2ZTGIf({
        \b6_2ZTGIf[147] }));
    b8_1LbcQDr1_x_77_0 b8_1LbcgKxJ (.mdiclink_reg({mdiclink_reg[77]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[77]}), .b4_nUAi({
        b4_nUAi[233], b4_nUAi[232], b4_nUAi[231]}), .b6_2ZTGIf({
        \b6_2ZTGIf[77] }));
    b8_1LbcQDr1_x_137_0 b8_1LbcgKGJ (.mdiclink_reg({mdiclink_reg[17]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[137]}), .b4_nUAi({
        b4_nUAi[52], b4_nUAi[51]}), .N_27(N_27_6), .N_25(N_25_6));
    b8_1LbcQDr1_x_100_0 b8_1LbcgKIQ0 (.mdiclink_reg({mdiclink_reg[54]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[100]}), .b4_nUAi({
        b4_nUAi[164], b4_nUAi[163], b4_nUAi[162]}), .b6_2ZTGIf({
        \b6_2ZTGIf[54] }));
    b8_1LbcQDr1_x_152_0 b7_1LbcgKw (.mdiclink_reg({mdiclink_reg[2]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[152]}), .b4_nUAi({b4_nUAi[7], 
        b4_nUAi[6]}), .N_27(N_27_1), .N_25(N_25_1));
    b8_1LbcQDr1_x_97_0 b8_1LbcgKIJ (.mdiclink_reg({mdiclink_reg[57]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[97]}), .b4_nUAi({
        b4_nUAi[173], b4_nUAi[172], b4_nUAi[171]}), .b6_2ZTGIf({
        \b6_2ZTGIf[57] }));
    b8_1LbcQDr1_x_14_0 b9_1LbcgKGQm0 (.mdiclink_reg({mdiclink_reg[140]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[14]}), .b4_nUAi({
        b4_nUAi[422], b4_nUAi[421], b4_nUAi[420]}), .b6_2ZTGIf({
        \b6_2ZTGIf[140] }));
    b8_1LbcQDr1_x_116_0 b8_1LbcgKen (.mdiclink_reg({mdiclink_reg[38]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[116]}), .b4_nUAi({
        b4_nUAi[116], b4_nUAi[115], b4_nUAi[114]}), .b6_2ZTGIf({
        \b6_2ZTGIf[38] }));
    b8_1LbcQDr1_x_68_0 b8_1LbcgKbA (.mdiclink_reg({mdiclink_reg[86]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[68]}), .b4_nUAi({
        b4_nUAi[260], b4_nUAi[259], b4_nUAi[258]}), .b6_2ZTGIf({
        \b6_2ZTGIf[86] }));
    b8_1LbcQDr1_x_112_0 b8_1LbcgKEI0 (.mdiclink_reg({mdiclink_reg[42]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[112]}), .b4_nUAi({
        b4_nUAi[127], b4_nUAi[126]}), .N_27(N_27_16), .N_25(N_25_16));
    b8_1LbcQDr1_x_19_0 b9_1LbcgKGqp (.mdiclink_reg({mdiclink_reg[135]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[19]}), .b4_nUAi({
        b4_nUAi[407], b4_nUAi[406], b4_nUAi[405]}), .b6_2ZTGIf({
        \b6_2ZTGIf[135] }));
    b8_1LbcQDr1_x_115_0 b8_1LbcgKeV (.mdiclink_reg({mdiclink_reg[39]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[115]}), .b4_nUAi({
        b4_nUAi[119], b4_nUAi[118], b4_nUAi[117]}), .b6_2ZTGIf({
        \b6_2ZTGIf[39] }));
    b8_1LbcQDr1_x_13_0 b9_1LbcgKGQn0 (.mdiclink_reg({mdiclink_reg[141]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[13]}), .b4_nUAi({
        b4_nUAi[425], b4_nUAi[424], b4_nUAi[423]}), .b6_2ZTGIf({
        \b6_2ZTGIf[141] }));
    b8_1LbcQDr1_x_15_0 b9_1LbcgKGqq (.mdiclink_reg({mdiclink_reg[139]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[15]}), .b4_nUAi({
        b4_nUAi[419], b4_nUAi[418], b4_nUAi[417]}), .b6_2ZTGIf({
        \b6_2ZTGIf[139] }));
    b8_1LbcQDr1_x_42_0 b9_1LbcgKGSd (.mdiclink_reg({mdiclink_reg[112]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[42]}), .b4_nUAi({
        b4_nUAi[337], b4_nUAi[336]}), .N_27(N_27_41), .N_25(N_25_41));
    b8_1LbcQDr1_x_0_0 b9_1LbcgKGUl (.mdiclink_reg({mdiclink_reg[154]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[0]}), .b4_nUAi({b4_nUAi[463], 
        b4_nUAi[462]}), .b6_2ZTGIf({\b6_2ZTGIf[154] }), .b7_PSyi3wy(
        b7_PSyi3wy));
    b8_1LbcQDr1_x_52_0 b9_1LbcgKGRd (.mdiclink_reg({mdiclink_reg[102]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[52]}), .b4_nUAi({
        b4_nUAi[308], b4_nUAi[307], b4_nUAi[306]}), .b6_2ZTGIf({
        \b6_2ZTGIf[102] }));
    b8_1LbcQDr1_x_16_0 b9_1LbcgKGqS (.mdiclink_reg({mdiclink_reg[138]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[16]}), .b4_nUAi({
        b4_nUAi[415], b4_nUAi[414]}), .N_27(N_27_52), .N_25(N_25_52));
    b8_1LbcQDr1_x_17_0 b9_1LbcgKGqe (.mdiclink_reg({mdiclink_reg[137]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[17]}), .b4_nUAi({
        b4_nUAi[413], b4_nUAi[412], b4_nUAi[411]}), .b6_2ZTGIf({
        \b6_2ZTGIf[137] }));
    b8_1LbcQDr1_x_128_0 b8_1LbcgKwA (.mdiclink_reg({mdiclink_reg[26]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[128]}), .b4_nUAi({
        b4_nUAi[79], b4_nUAi[78]}), .N_27(N_27_10), .N_25(N_25_10));
    b8_1LbcQDr1_x_154_0 b7_1LbcgKF (.mdiclink_reg({mdiclink_reg[0]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[154]}), .b4_nUAi({b4_nUAi[1], 
        b4_nUAi[0]}), .N_27(N_27), .N_25(N_25));
    b8_1LbcQDr1_x_24_0 b9_1LbcgKGqm (.mdiclink_reg({mdiclink_reg[130]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[24]}), .b4_nUAi({
        b4_nUAi[391], b4_nUAi[390]}), .N_27(N_27_49), .N_25(N_25_49));
    b8_1LbcQDr1_x_88_0 b8_1LbcgKoA (.mdiclink_reg({mdiclink_reg[66]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[88]}), .b4_nUAi({
        b4_nUAi[199], b4_nUAi[198]}), .N_27(N_27_25), .N_25(N_25_25));
    b8_1LbcQDr1_x_39_0 b9_1LbcgKGSp (.mdiclink_reg({mdiclink_reg[115]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[39]}), .b4_nUAi({
        b4_nUAi[346], b4_nUAi[345]}), .N_27(N_27_44), .N_25(N_25_44));
    b8_1LbcQDr1_x_49_0 b9_1LbcgKGRp (.mdiclink_reg({mdiclink_reg[105]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[49]}), .b4_nUAi({
        b4_nUAi[317], b4_nUAi[316], b4_nUAi[315]}), .b6_2ZTGIf({
        \b6_2ZTGIf[105] }));
    b8_1LbcQDr1_x_56_0 b8_1LbcgKJn (.mdiclink_reg({mdiclink_reg[98]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[56]}), .b4_nUAi({
        b4_nUAi[295], b4_nUAi[294]}), .N_27(N_27_37), .N_25(N_25_37));
    b8_1LbcQDr1_x_71_0 b8_1LbcgKbq (.mdiclink_reg({mdiclink_reg[83]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[71]}), .b4_nUAi({
        b4_nUAi[250], b4_nUAi[249]}), .N_27(N_27_32), .N_25(N_25_32));
    b8_1LbcQDr1_x_30_0 b9_1LbcgKGIl (.mdiclink_reg({mdiclink_reg[124]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[30]}), .b4_nUAi({
        b4_nUAi[374], b4_nUAi[373], b4_nUAi[372]}), .b6_2ZTGIf({
        \b6_2ZTGIf[124] }));
    b8_1LbcQDr1_x_107_0 b8_1LbcgKEJ0 (.mdiclink_reg({mdiclink_reg[47]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[107]}), .b4_nUAi({
        b4_nUAi[143], b4_nUAi[142], b4_nUAi[141]}), .b6_2ZTGIf({
        \b6_2ZTGIf[47] }));
    b8_1LbcQDr1_x_35_0 b9_1LbcgKGSq (.mdiclink_reg({mdiclink_reg[119]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[35]}), .b4_nUAi({
        b4_nUAi[359], b4_nUAi[358], b4_nUAi[357]}), .b6_2ZTGIf({
        \b6_2ZTGIf[119] }));
    b8_1LbcQDr1_x_28_0 b9_1LbcgKGI5 (.mdiclink_reg({mdiclink_reg[126]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[28]}), .b4_nUAi({
        b4_nUAi[380], b4_nUAi[379], b4_nUAi[378]}), .b6_2ZTGIf({
        \b6_2ZTGIf[126] }));
    b8_1LbcQDr1_x_23_0 b9_1LbcgKGqn (.mdiclink_reg({mdiclink_reg[131]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[23]}), .b4_nUAi({
        b4_nUAi[394], b4_nUAi[393]}), .N_27(N_27_50), .N_25(N_25_50));
    b8_1LbcQDr1_x_45_0 b9_1LbcgKGRq (.mdiclink_reg({mdiclink_reg[109]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[45]}), .b4_nUAi({
        b4_nUAi[329], b4_nUAi[328], b4_nUAi[327]}), .b6_2ZTGIf({
        \b6_2ZTGIf[109] }));
    b8_1LbcQDr1_x_36_0 b9_1LbcgKGSS (.mdiclink_reg({mdiclink_reg[118]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[36]}), .b4_nUAi({
        b4_nUAi[356], b4_nUAi[355], b4_nUAi[354]}), .b6_2ZTGIf({
        \b6_2ZTGIf[118] }));
    b8_1LbcQDr1_x_55_0 b8_1LbcgKJV (.mdiclink_reg({mdiclink_reg[99]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[55]}), .b4_nUAi({
        b4_nUAi[298], b4_nUAi[297]}), .N_27(N_27_38), .N_25(N_25_38));
    b8_1LbcQDr1_x_119_0 b8_1LbcgKeU (.mdiclink_reg({mdiclink_reg[35]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[119]}), .b4_nUAi({
        b4_nUAi[106], b4_nUAi[105]}), .N_27(N_27_14), .N_25(N_25_14));
    b8_1LbcQDr1_x_46_0 b9_1LbcgKGRS (.mdiclink_reg({mdiclink_reg[108]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[46]}), .b4_nUAi({
        b4_nUAi[326], b4_nUAi[325], b4_nUAi[324]}), .b6_2ZTGIf({
        \b6_2ZTGIf[108] }));
    b8_1LbcQDr1_x_151_0 b7_1LbcgKe (.mdiclink_reg({mdiclink_reg[3]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[151]}), .b4_nUAi({
        b4_nUAi[10], b4_nUAi[9]}), .N_27(N_27_2), .N_25(N_25_2));
    b8_1LbcQDr1_x_37_0 b9_1LbcgKGSe (.mdiclink_reg({mdiclink_reg[117]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[37]}), .b4_nUAi({
        b4_nUAi[353], b4_nUAi[352], b4_nUAi[351]}), .b6_2ZTGIf({
        \b6_2ZTGIf[117] }));
    b8_1LbcQDr1_x_11_0 b9_1LbcgKGQV0 (.mdiclink_reg({mdiclink_reg[143]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[11]}), .b4_nUAi({
        b4_nUAi[431], b4_nUAi[430], b4_nUAi[429]}), .b6_2ZTGIf({
        \b6_2ZTGIf[143] }));
    b8_1LbcQDr1_x_47_0 b9_1LbcgKGRe (.mdiclink_reg({mdiclink_reg[107]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[47]}), .b4_nUAi({
        b4_nUAi[323], b4_nUAi[322], b4_nUAi[321]}), .b6_2ZTGIf({
        \b6_2ZTGIf[107] }));
    b8_1LbcQDr1_x_44_0 b9_1LbcgKGSm (.mdiclink_reg({mdiclink_reg[110]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[44]}), .b4_nUAi({
        b4_nUAi[332], b4_nUAi[331], b4_nUAi[330]}), .b6_2ZTGIf({
        \b6_2ZTGIf[110] }));
    b8_1LbcQDr1_x_54_0 b9_1LbcgKGRm (.mdiclink_reg({mdiclink_reg[100]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[54]}), .b4_nUAi({
        b4_nUAi[302], b4_nUAi[301], b4_nUAi[300]}), .b6_2ZTGIf({
        \b6_2ZTGIf[100] }));
    b8_1LbcQDr1_x_73_0 b8_1LbcgKbS (.mdiclink_reg({mdiclink_reg[81]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[73]}), .b4_nUAi({
        b4_nUAi[244], b4_nUAi[243]}), .N_27(N_27_30), .N_25(N_25_30));
    b8_1LbcQDr1_x_74_0 b8_1LbcgKbR (.mdiclink_reg({mdiclink_reg[80]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[74]}), .b4_nUAi({
        b4_nUAi[241], b4_nUAi[240]}), .N_27(N_27_29), .N_25(N_25_29));
    b8_1LbcQDr1_x_122_0 b8_1LbcgKeI (.mdiclink_reg({mdiclink_reg[32]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[122]}), .b4_nUAi({
        b4_nUAi[97], b4_nUAi[96]}), .N_27(N_27_11), .N_25(N_25_11));
    b8_1LbcQDr1_x_43_0 b9_1LbcgKGSn (.mdiclink_reg({mdiclink_reg[111]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[43]}), .b4_nUAi({
        b4_nUAi[335], b4_nUAi[334], b4_nUAi[333]}), .b6_2ZTGIf({
        \b6_2ZTGIf[111] }));
    b8_1LbcQDr1_x_131_0 b8_1LbcgKwq (.mdiclink_reg({mdiclink_reg[23]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[131]}), .b4_nUAi({
        b4_nUAi[71], b4_nUAi[70], b4_nUAi[69]}), .b6_2ZTGIf({
        \b6_2ZTGIf[23] }));
    b8_1LbcQDr1_x_91_0 b8_1LbcgKoq (.mdiclink_reg({mdiclink_reg[63]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[91]}), .b4_nUAi({
        b4_nUAi[191], b4_nUAi[190], b4_nUAi[189]}), .b6_2ZTGIf({
        \b6_2ZTGIf[63] }));
    b8_1LbcQDr1_x_53_0 b9_1LbcgKGRn (.mdiclink_reg({mdiclink_reg[101]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[53]}), .b4_nUAi({
        b4_nUAi[305], b4_nUAi[304], b4_nUAi[303]}), .b6_2ZTGIf({
        \b6_2ZTGIf[101] }));
    b8_1LbcQDr1_x_21_0 b9_1LbcgKGqV (.mdiclink_reg({mdiclink_reg[133]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[21]}), .b4_nUAi({
        b4_nUAi[401], b4_nUAi[400], b4_nUAi[399]}), .b6_2ZTGIf({
        \b6_2ZTGIf[133] }));
    b8_1LbcQDr1_x_59_0 b8_1LbcgKJU (.mdiclink_reg({mdiclink_reg[95]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[59]}), .b4_nUAi({
        b4_nUAi[287], b4_nUAi[286], b4_nUAi[285]}), .b6_2ZTGIf({
        \b6_2ZTGIf[95] }));
    b8_1LbcQDr1_x_146_0 b7_1LbcgKb (.mdiclink_reg({mdiclink_reg[8]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[146]}), .b4_nUAi({
        b4_nUAi[25], b4_nUAi[24]}), .N_27(N_27_3), .N_25(N_25_3));
    b8_1LbcQDr1_x_133_0 b8_1LbcgKwS (.mdiclink_reg({mdiclink_reg[21]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[133]}), .b4_nUAi({
        b4_nUAi[65], b4_nUAi[64], b4_nUAi[63]}), .b6_2ZTGIf({
        \b6_2ZTGIf[21] }));
    b8_1LbcQDr1_x_93_0 b8_1LbcgKoS (.mdiclink_reg({mdiclink_reg[61]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[93]}), .b4_nUAi({
        b4_nUAi[185], b4_nUAi[184], b4_nUAi[183]}), .b6_2ZTGIf({
        \b6_2ZTGIf[61] }));
    b8_1LbcQDr1_x_134_0 b8_1LbcgKwR (.mdiclink_reg({mdiclink_reg[20]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[134]}), .b4_nUAi({
        b4_nUAi[62], b4_nUAi[61], b4_nUAi[60]}), .b6_2ZTGIf({
        \b6_2ZTGIf[20] }));
    b8_1LbcQDr1_x_94_0 b8_1LbcgKoR (.mdiclink_reg({mdiclink_reg[60]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[94]}), .b4_nUAi({
        b4_nUAi[182], b4_nUAi[181], b4_nUAi[180]}), .b6_2ZTGIf({
        \b6_2ZTGIf[60] }));
    b8_1LbcQDr1_x_62_0 b8_1LbcgKJI (.mdiclink_reg({mdiclink_reg[92]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[62]}), .b4_nUAi({
        b4_nUAi[278], b4_nUAi[277], b4_nUAi[276]}), .b6_2ZTGIf({
        \b6_2ZTGIf[92] }));
    b8_1LbcQDr1_x_78_0 b8_1LbcgKxA (.mdiclink_reg({mdiclink_reg[76]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[78]}), .b4_nUAi({
        b4_nUAi[230], b4_nUAi[229], b4_nUAi[228]}), .b6_2ZTGIf({
        \b6_2ZTGIf[76] }));
    b8_1LbcQDr1_x_138_0 b8_1LbcgKGA (.mdiclink_reg({mdiclink_reg[16]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[138]}), .b4_nUAi({
        b4_nUAi[49], b4_nUAi[48]}), .N_27(N_27_5), .N_25(N_25_5));
    b8_1LbcQDr1_x_117_0 b8_1LbcgKeJ (.mdiclink_reg({mdiclink_reg[37]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[117]}), .b4_nUAi({
        b4_nUAi[113], b4_nUAi[112], b4_nUAi[111]}), .b6_2ZTGIf({
        \b6_2ZTGIf[37] }));
    b8_1LbcQDr1_x_41_0 b9_1LbcgKGSV (.mdiclink_reg({mdiclink_reg[113]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[41]}), .b4_nUAi({
        b4_nUAi[340], b4_nUAi[339]}), .N_27(N_27_42), .N_25(N_25_42));
    b8_1LbcQDr1_x_66_0 b8_1LbcgKbn (.mdiclink_reg({mdiclink_reg[88]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[66]}), .b4_nUAi({
        b4_nUAi[265], b4_nUAi[264]}), .N_27(N_27_33), .N_25(N_25_33));
    b8_1LbcQDr1_x_51_0 b9_1LbcgKGRV (.mdiclink_reg({mdiclink_reg[103]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[51]}), .b4_nUAi({
        b4_nUAi[311], b4_nUAi[310], b4_nUAi[309]}), .b6_2ZTGIf({
        \b6_2ZTGIf[103] }));
    b8_1LbcQDr1_x_98_0 b8_1LbcgKIA (.mdiclink_reg({mdiclink_reg[56]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[98]}), .b4_nUAi({
        b4_nUAi[169], b4_nUAi[168]}), .N_27(N_27_21), .N_25(N_25_21));
    b8_1LbcQDr1_x_70_0 b8_1LbcgKbQ0 (.mdiclink_reg({mdiclink_reg[84]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[70]}), .b4_nUAi({
        b4_nUAi[254], b4_nUAi[253], b4_nUAi[252]}), .b6_2ZTGIf({
        \b6_2ZTGIf[84] }));
    b8_1LbcQDr1_x_2_0 b9_1LbcgKGUd (.mdiclink_reg({mdiclink_reg[152]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[2]}), .b4_nUAi({b4_nUAi[458], 
        b4_nUAi[457], b4_nUAi[456]}), .b6_2ZTGIf({\b6_2ZTGIf[152] }));
    b8_1LbcQDr1_x_65_0 b8_1LbcgKbV (.mdiclink_reg({mdiclink_reg[89]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[65]}), .b4_nUAi({
        b4_nUAi[269], b4_nUAi[268], b4_nUAi[267]}), .b6_2ZTGIf({
        \b6_2ZTGIf[89] }));
    b8_1LbcQDr1_x_153_0 b7_1LbcgKG (.mdiclink_reg({mdiclink_reg[1]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[153]}), .b4_nUAi({b4_nUAi[4], 
        b4_nUAi[3]}), .N_27(N_27_0), .N_25(N_25_0));
    b8_1LbcQDr1_x_60_0 b8_1LbcgKJQ0 (.mdiclink_reg({mdiclink_reg[94]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[60]}), .b4_nUAi({
        b4_nUAi[284], b4_nUAi[283], b4_nUAi[282]}), .b6_2ZTGIf({
        \b6_2ZTGIf[94] }));
    b8_1LbcQDr1_x_32_0 b9_1LbcgKGId (.mdiclink_reg({mdiclink_reg[122]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[32]}), .b4_nUAi({
        b4_nUAi[367], b4_nUAi[366]}), .N_27(N_27_46), .N_25(N_25_46));
    b8_1LbcQDr1_x_145_0 b7_1LbcgKJ (.mdiclink_reg({mdiclink_reg[9]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[145]}), .b4_nUAi({
        b4_nUAi[29], b4_nUAi[28], b4_nUAi[27]}), .b6_2ZTGIf({
        \b6_2ZTGIf[9] }));
    b8_1LbcQDr1_x_126_0 b8_1LbcgKwn (.mdiclink_reg({mdiclink_reg[28]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[126]}), .b4_nUAi({
        b4_nUAi[86], b4_nUAi[85], b4_nUAi[84]}), .b6_2ZTGIf({
        \b6_2ZTGIf[28] }));
    b8_1LbcQDr1_x_86_0 b8_1LbcgKon (.mdiclink_reg({mdiclink_reg[68]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[86]}), .b4_nUAi({
        b4_nUAi[206], b4_nUAi[205], b4_nUAi[204]}), .b6_2ZTGIf({
        \b6_2ZTGIf[68] }));
    b8_1LbcQDr1_x_57_0 b8_1LbcgKJJ (.mdiclink_reg({mdiclink_reg[97]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[57]}), .b4_nUAi({
        b4_nUAi[292], b4_nUAi[291]}), .N_27(N_27_36), .N_25(N_25_36));
    b8_1LbcQDr1_x_81_0 b8_1LbcgKxq (.mdiclink_reg({mdiclink_reg[73]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[81]}), .b4_nUAi({
        b4_nUAi[221], b4_nUAi[220], b4_nUAi[219]}), .b6_2ZTGIf({
        \b6_2ZTGIf[73] }));
    b8_1LbcQDr1_x_141_0 b8_1LbcgKGq (.mdiclink_reg({mdiclink_reg[13]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[141]}), .b4_nUAi({
        b4_nUAi[41], b4_nUAi[40], b4_nUAi[39]}), .b6_2ZTGIf({
        \b6_2ZTGIf[13] }));
    b8_1LbcQDr1_x_111_0 b8_1LbcgKEq0 (.mdiclink_reg({mdiclink_reg[43]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[111]}), .b4_nUAi({
        b4_nUAi[131], b4_nUAi[130], b4_nUAi[129]}), .b6_2ZTGIf({
        \b6_2ZTGIf[43] }));
    b8_1LbcQDr1_x_29_0 b9_1LbcgKGIp (.mdiclink_reg({mdiclink_reg[125]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[29]}), .b4_nUAi({
        b4_nUAi[377], b4_nUAi[376], b4_nUAi[375]}), .b6_2ZTGIf({
        \b6_2ZTGIf[125] }));
    b8_1LbcQDr1_x_101_0 b8_1LbcgKIq (.mdiclink_reg({mdiclink_reg[53]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[101]}), .b4_nUAi({
        b4_nUAi[161], b4_nUAi[160], b4_nUAi[159]}), .b6_2ZTGIf({
        \b6_2ZTGIf[53] }));
    b8_1LbcQDr1_x_125_0 b8_1LbcgKwV (.mdiclink_reg({mdiclink_reg[29]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[125]}), .b4_nUAi({
        b4_nUAi[89], b4_nUAi[88], b4_nUAi[87]}), .b6_2ZTGIf({
        \b6_2ZTGIf[29] }));
    b8_1LbcQDr1_x_4_0 b9_1LbcgKGUm (.mdiclink_reg({mdiclink_reg[150]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[4]}), .b4_nUAi({b4_nUAi[451], 
        b4_nUAi[450]}), .N_27(N_27_55), .N_25(N_25_55));
    b8_1LbcQDr1_x_85_0 b8_1LbcgKoV (.mdiclink_reg({mdiclink_reg[69]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[85]}), .b4_nUAi({
        b4_nUAi[209], b4_nUAi[208], b4_nUAi[207]}), .b6_2ZTGIf({
        \b6_2ZTGIf[69] }));
    b8_1LbcQDr1_x_108_0 b8_1LbcgKEA0 (.mdiclink_reg({mdiclink_reg[46]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[108]}), .b4_nUAi({
        b4_nUAi[140], b4_nUAi[139], b4_nUAi[138]}), .b6_2ZTGIf({
        \b6_2ZTGIf[46] }));
    b8_1LbcQDr1_x_25_0 b9_1LbcgKGIq (.mdiclink_reg({mdiclink_reg[129]})
        , .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[25]}), .b4_nUAi({
        b4_nUAi[388], b4_nUAi[387]}), .N_27(N_27_48), .N_25(N_25_48));
    b8_1LbcQDr1_x_69_0 b8_1LbcgKbU (.mdiclink_reg({mdiclink_reg[85]}), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[69]}), .b4_nUAi({
        b4_nUAi[257], b4_nUAi[256], b4_nUAi[255]}), .b6_2ZTGIf({
        \b6_2ZTGIf[85] }));
    
endmodule


module b7_PfFzrNY_x_0(
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       IICE_comm2iice,
       b11_PSyil9s_FMZ,
       BW_clk_c,
       b7_PSyi3wy,
       b4_PLyF,
       b8_PSyiBgYG
    );
input  [154:0] mdiclink_reg;
input  [154:0] b11_OFWNT9L_8tZ;
input  [11:10] IICE_comm2iice;
output b11_PSyil9s_FMZ;
input  BW_clk_c;
output b7_PSyi3wy;
input  b4_PLyF;
input  b8_PSyiBgYG;

    wire VCC_net_1, \b11_uUT0JC4gFrY[1] , GND_net_1, \b4_nUAi[0] , 
        \b4_nUAi[1] , \b4_nUAi[2] , \b4_nUAi[3] , \b4_nUAi[4] , 
        \b4_nUAi[5] , \b4_nUAi[6] , \b4_nUAi[7] , \b4_nUAi[8] , 
        \b4_nUAi[9] , \b4_nUAi[10] , \b4_nUAi[11] , \b4_nUAi[12] , 
        \b4_nUAi[13] , \b4_nUAi[14] , \b4_nUAi[15] , \b4_nUAi[16] , 
        \b4_nUAi[17] , \b4_nUAi[18] , \b4_nUAi[19] , \b4_nUAi[20] , 
        \b4_nUAi[21] , \b4_nUAi[22] , \b4_nUAi[23] , \b4_nUAi[24] , 
        \b4_nUAi[25] , \b4_nUAi[26] , \b4_nUAi[27] , \b4_nUAi[28] , 
        \b4_nUAi[29] , \b4_nUAi[30] , \b4_nUAi[31] , \b4_nUAi[32] , 
        \b4_nUAi[33] , \b4_nUAi[34] , \b4_nUAi[35] , \b4_nUAi[36] , 
        \b4_nUAi[37] , \b4_nUAi[38] , \b4_nUAi[39] , \b4_nUAi[40] , 
        \b4_nUAi[41] , \b4_nUAi[42] , \b4_nUAi[43] , \b4_nUAi[44] , 
        \b4_nUAi[45] , \b4_nUAi[46] , \b4_nUAi[47] , \b4_nUAi[48] , 
        \b4_nUAi[49] , \b4_nUAi[50] , \b4_nUAi[51] , \b4_nUAi[52] , 
        \b4_nUAi[53] , \b4_nUAi[54] , \b4_nUAi[55] , \b4_nUAi[56] , 
        \b4_nUAi[57] , \b4_nUAi[58] , \b4_nUAi[59] , \b4_nUAi[60] , 
        \b4_nUAi[61] , \b4_nUAi[62] , \b4_nUAi[63] , \b4_nUAi[64] , 
        \b4_nUAi[65] , \b4_nUAi[66] , \b4_nUAi[67] , \b4_nUAi[68] , 
        \b4_nUAi[69] , \b4_nUAi[70] , \b4_nUAi[71] , \b4_nUAi[72] , 
        \b4_nUAi[73] , \b4_nUAi[74] , \b4_nUAi[75] , \b4_nUAi[76] , 
        \b4_nUAi[77] , \b4_nUAi[78] , \b4_nUAi[79] , \b4_nUAi[80] , 
        \b4_nUAi[81] , \b4_nUAi[82] , \b4_nUAi[83] , \b4_nUAi[84] , 
        \b4_nUAi[85] , \b4_nUAi[86] , \b4_nUAi[87] , \b4_nUAi[88] , 
        \b4_nUAi[89] , \b4_nUAi[90] , \b4_nUAi[91] , \b4_nUAi[92] , 
        \b4_nUAi[93] , \b4_nUAi[94] , \b4_nUAi[95] , \b4_nUAi[96] , 
        \b4_nUAi[97] , \b4_nUAi[98] , \b4_nUAi[99] , \b4_nUAi[100] , 
        \b4_nUAi[101] , \b4_nUAi[102] , \b4_nUAi[103] , \b4_nUAi[104] , 
        \b4_nUAi[105] , \b4_nUAi[106] , \b4_nUAi[107] , \b4_nUAi[108] , 
        \b4_nUAi[109] , \b4_nUAi[110] , \b4_nUAi[111] , \b4_nUAi[112] , 
        \b4_nUAi[113] , \b4_nUAi[114] , \b4_nUAi[115] , \b4_nUAi[116] , 
        \b4_nUAi[117] , \b4_nUAi[118] , \b4_nUAi[119] , \b4_nUAi[120] , 
        \b4_nUAi[121] , \b4_nUAi[122] , \b4_nUAi[123] , \b4_nUAi[124] , 
        \b4_nUAi[125] , \b4_nUAi[126] , \b4_nUAi[127] , \b4_nUAi[128] , 
        \b4_nUAi[129] , \b4_nUAi[130] , \b4_nUAi[131] , \b4_nUAi[132] , 
        \b4_nUAi[133] , \b4_nUAi[134] , \b4_nUAi[135] , \b4_nUAi[136] , 
        \b4_nUAi[137] , \b4_nUAi[138] , \b4_nUAi[139] , \b4_nUAi[140] , 
        \b4_nUAi[141] , \b4_nUAi[142] , \b4_nUAi[143] , \b4_nUAi[144] , 
        \b4_nUAi[145] , \b4_nUAi[146] , \b4_nUAi[147] , \b4_nUAi[148] , 
        \b4_nUAi[149] , \b4_nUAi[150] , \b4_nUAi[151] , \b4_nUAi[152] , 
        \b4_nUAi[153] , \b4_nUAi[154] , \b4_nUAi[155] , \b4_nUAi[156] , 
        \b4_nUAi[157] , \b4_nUAi[158] , \b4_nUAi[159] , \b4_nUAi[160] , 
        \b4_nUAi[161] , \b4_nUAi[162] , \b4_nUAi[163] , \b4_nUAi[164] , 
        \b4_nUAi[165] , \b4_nUAi[166] , \b4_nUAi[167] , \b4_nUAi[168] , 
        \b4_nUAi[169] , \b4_nUAi[170] , \b4_nUAi[171] , \b4_nUAi[172] , 
        \b4_nUAi[173] , \b4_nUAi[174] , \b4_nUAi[175] , \b4_nUAi[176] , 
        \b4_nUAi[177] , \b4_nUAi[178] , \b4_nUAi[179] , \b4_nUAi[180] , 
        \b4_nUAi[181] , \b4_nUAi[182] , \b4_nUAi[183] , \b4_nUAi[184] , 
        \b4_nUAi[185] , \b4_nUAi[186] , \b4_nUAi[187] , \b4_nUAi[188] , 
        \b4_nUAi[189] , \b4_nUAi[190] , \b4_nUAi[191] , \b4_nUAi[192] , 
        \b4_nUAi[193] , \b4_nUAi[194] , \b4_nUAi[195] , \b4_nUAi[196] , 
        \b4_nUAi[197] , \b4_nUAi[198] , \b4_nUAi[199] , \b4_nUAi[200] , 
        \b4_nUAi[201] , \b4_nUAi[202] , \b4_nUAi[203] , \b4_nUAi[204] , 
        \b4_nUAi[205] , \b4_nUAi[206] , \b4_nUAi[207] , \b4_nUAi[208] , 
        \b4_nUAi[209] , \b4_nUAi[210] , \b4_nUAi[211] , \b4_nUAi[212] , 
        \b4_nUAi[213] , \b4_nUAi[214] , \b4_nUAi[215] , \b4_nUAi[216] , 
        \b4_nUAi[217] , \b4_nUAi[218] , \b4_nUAi[219] , \b4_nUAi[220] , 
        \b4_nUAi[221] , \b4_nUAi[222] , \b4_nUAi[223] , \b4_nUAi[224] , 
        \b4_nUAi[225] , \b4_nUAi[226] , \b4_nUAi[227] , \b4_nUAi[228] , 
        \b4_nUAi[229] , \b4_nUAi[230] , \b4_nUAi[231] , \b4_nUAi[232] , 
        \b4_nUAi[233] , \b4_nUAi[234] , \b4_nUAi[235] , \b4_nUAi[236] , 
        \b4_nUAi[237] , \b4_nUAi[238] , \b4_nUAi[239] , \b4_nUAi[240] , 
        \b4_nUAi[241] , \b4_nUAi[242] , \b4_nUAi[243] , \b4_nUAi[244] , 
        \b4_nUAi[245] , \b4_nUAi[246] , \b4_nUAi[247] , \b4_nUAi[248] , 
        \b4_nUAi[249] , \b4_nUAi[250] , \b4_nUAi[251] , \b4_nUAi[252] , 
        \b4_nUAi[253] , \b4_nUAi[254] , \b4_nUAi[255] , \b4_nUAi[256] , 
        \b4_nUAi[257] , \b4_nUAi[258] , \b4_nUAi[259] , \b4_nUAi[260] , 
        \b4_nUAi[261] , \b4_nUAi[262] , \b4_nUAi[263] , \b4_nUAi[264] , 
        \b4_nUAi[265] , \b4_nUAi[266] , \b4_nUAi[267] , \b4_nUAi[268] , 
        \b4_nUAi[269] , \b4_nUAi[270] , \b4_nUAi[271] , \b4_nUAi[272] , 
        \b4_nUAi[273] , \b4_nUAi[274] , \b4_nUAi[275] , \b4_nUAi[276] , 
        \b4_nUAi[277] , \b4_nUAi[278] , \b4_nUAi[279] , \b4_nUAi[280] , 
        \b4_nUAi[281] , \b4_nUAi[282] , \b4_nUAi[283] , \b4_nUAi[284] , 
        \b4_nUAi[285] , \b4_nUAi[286] , \b4_nUAi[287] , \b4_nUAi[288] , 
        \b4_nUAi[289] , \b4_nUAi[290] , \b4_nUAi[291] , \b4_nUAi[292] , 
        \b4_nUAi[293] , \b4_nUAi[294] , \b4_nUAi[295] , \b4_nUAi[296] , 
        \b4_nUAi[297] , \b4_nUAi[298] , \b4_nUAi[299] , \b4_nUAi[300] , 
        \b4_nUAi[301] , \b4_nUAi[302] , \b4_nUAi[303] , \b4_nUAi[304] , 
        \b4_nUAi[305] , \b4_nUAi[306] , \b4_nUAi[307] , \b4_nUAi[308] , 
        \b4_nUAi[309] , \b4_nUAi[310] , \b4_nUAi[311] , \b4_nUAi[312] , 
        \b4_nUAi[313] , \b4_nUAi[314] , \b4_nUAi[315] , \b4_nUAi[316] , 
        \b4_nUAi[317] , \b4_nUAi[318] , \b4_nUAi[319] , \b4_nUAi[320] , 
        \b4_nUAi[321] , \b4_nUAi[322] , \b4_nUAi[323] , \b4_nUAi[324] , 
        \b4_nUAi[325] , \b4_nUAi[326] , \b4_nUAi[327] , \b4_nUAi[328] , 
        \b4_nUAi[329] , \b4_nUAi[330] , \b4_nUAi[331] , \b4_nUAi[332] , 
        \b4_nUAi[333] , \b4_nUAi[334] , \b4_nUAi[335] , \b4_nUAi[336] , 
        \b4_nUAi[337] , \b4_nUAi[338] , \b4_nUAi[339] , \b4_nUAi[340] , 
        \b4_nUAi[341] , \b4_nUAi[342] , \b4_nUAi[343] , \b4_nUAi[344] , 
        \b4_nUAi[345] , \b4_nUAi[346] , \b4_nUAi[347] , \b4_nUAi[348] , 
        \b4_nUAi[349] , \b4_nUAi[350] , \b4_nUAi[351] , \b4_nUAi[352] , 
        \b4_nUAi[353] , \b4_nUAi[354] , \b4_nUAi[355] , \b4_nUAi[356] , 
        \b4_nUAi[357] , \b4_nUAi[358] , \b4_nUAi[359] , \b4_nUAi[360] , 
        \b4_nUAi[361] , \b4_nUAi[362] , \b4_nUAi[363] , \b4_nUAi[364] , 
        \b4_nUAi[365] , \b4_nUAi[366] , \b4_nUAi[367] , \b4_nUAi[368] , 
        \b4_nUAi[369] , \b4_nUAi[370] , \b4_nUAi[371] , \b4_nUAi[372] , 
        \b4_nUAi[373] , \b4_nUAi[374] , \b4_nUAi[375] , \b4_nUAi[376] , 
        \b4_nUAi[377] , \b4_nUAi[378] , \b4_nUAi[379] , \b4_nUAi[380] , 
        \b4_nUAi[381] , \b4_nUAi[382] , \b4_nUAi[383] , \b4_nUAi[384] , 
        \b4_nUAi[385] , \b4_nUAi[386] , \b4_nUAi[387] , \b4_nUAi[388] , 
        \b4_nUAi[389] , \b4_nUAi[390] , \b4_nUAi[391] , \b4_nUAi[392] , 
        \b4_nUAi[393] , \b4_nUAi[394] , \b4_nUAi[395] , \b4_nUAi[396] , 
        \b4_nUAi[397] , \b4_nUAi[398] , \b4_nUAi[399] , \b4_nUAi[400] , 
        \b4_nUAi[401] , \b4_nUAi[402] , \b4_nUAi[403] , \b4_nUAi[404] , 
        \b4_nUAi[405] , \b4_nUAi[406] , \b4_nUAi[407] , \b4_nUAi[408] , 
        \b4_nUAi[409] , \b4_nUAi[410] , \b4_nUAi[411] , \b4_nUAi[412] , 
        \b4_nUAi[413] , \b4_nUAi[414] , \b4_nUAi[415] , \b4_nUAi[416] , 
        \b4_nUAi[417] , \b4_nUAi[418] , \b4_nUAi[419] , \b4_nUAi[420] , 
        \b4_nUAi[421] , \b4_nUAi[422] , \b4_nUAi[423] , \b4_nUAi[424] , 
        \b4_nUAi[425] , \b4_nUAi[426] , \b4_nUAi[427] , \b4_nUAi[428] , 
        \b4_nUAi[429] , \b4_nUAi[430] , \b4_nUAi[431] , \b4_nUAi[432] , 
        \b4_nUAi[433] , \b4_nUAi[434] , \b4_nUAi[435] , \b4_nUAi[436] , 
        \b4_nUAi[437] , \b4_nUAi[438] , \b4_nUAi[439] , \b4_nUAi[440] , 
        \b4_nUAi[441] , \b4_nUAi[442] , \b4_nUAi[443] , \b4_nUAi[444] , 
        \b4_nUAi[445] , \b4_nUAi[446] , \b4_nUAi[447] , \b4_nUAi[448] , 
        \b4_nUAi[449] , \b4_nUAi[450] , \b4_nUAi[451] , \b4_nUAi[452] , 
        \b4_nUAi[453] , \b4_nUAi[454] , \b4_nUAi[455] , \b4_nUAi[456] , 
        \b4_nUAi[457] , \b4_nUAi[458] , \b4_nUAi[459] , \b4_nUAi[460] , 
        \b4_nUAi[461] , \b4_nUAi[462] , \b4_nUAi[463] ;
    
    b5_nvmFL_465s_x_0 b5_PbrtL (.b4_nUAi({\b4_nUAi[463] , 
        \b4_nUAi[462] , \b4_nUAi[461] , \b4_nUAi[460] , \b4_nUAi[459] , 
        \b4_nUAi[458] , \b4_nUAi[457] , \b4_nUAi[456] , \b4_nUAi[455] , 
        \b4_nUAi[454] , \b4_nUAi[453] , \b4_nUAi[452] , \b4_nUAi[451] , 
        \b4_nUAi[450] , \b4_nUAi[449] , \b4_nUAi[448] , \b4_nUAi[447] , 
        \b4_nUAi[446] , \b4_nUAi[445] , \b4_nUAi[444] , \b4_nUAi[443] , 
        \b4_nUAi[442] , \b4_nUAi[441] , \b4_nUAi[440] , \b4_nUAi[439] , 
        \b4_nUAi[438] , \b4_nUAi[437] , \b4_nUAi[436] , \b4_nUAi[435] , 
        \b4_nUAi[434] , \b4_nUAi[433] , \b4_nUAi[432] , \b4_nUAi[431] , 
        \b4_nUAi[430] , \b4_nUAi[429] , \b4_nUAi[428] , \b4_nUAi[427] , 
        \b4_nUAi[426] , \b4_nUAi[425] , \b4_nUAi[424] , \b4_nUAi[423] , 
        \b4_nUAi[422] , \b4_nUAi[421] , \b4_nUAi[420] , \b4_nUAi[419] , 
        \b4_nUAi[418] , \b4_nUAi[417] , \b4_nUAi[416] , \b4_nUAi[415] , 
        \b4_nUAi[414] , \b4_nUAi[413] , \b4_nUAi[412] , \b4_nUAi[411] , 
        \b4_nUAi[410] , \b4_nUAi[409] , \b4_nUAi[408] , \b4_nUAi[407] , 
        \b4_nUAi[406] , \b4_nUAi[405] , \b4_nUAi[404] , \b4_nUAi[403] , 
        \b4_nUAi[402] , \b4_nUAi[401] , \b4_nUAi[400] , \b4_nUAi[399] , 
        \b4_nUAi[398] , \b4_nUAi[397] , \b4_nUAi[396] , \b4_nUAi[395] , 
        \b4_nUAi[394] , \b4_nUAi[393] , \b4_nUAi[392] , \b4_nUAi[391] , 
        \b4_nUAi[390] , \b4_nUAi[389] , \b4_nUAi[388] , \b4_nUAi[387] , 
        \b4_nUAi[386] , \b4_nUAi[385] , \b4_nUAi[384] , \b4_nUAi[383] , 
        \b4_nUAi[382] , \b4_nUAi[381] , \b4_nUAi[380] , \b4_nUAi[379] , 
        \b4_nUAi[378] , \b4_nUAi[377] , \b4_nUAi[376] , \b4_nUAi[375] , 
        \b4_nUAi[374] , \b4_nUAi[373] , \b4_nUAi[372] , \b4_nUAi[371] , 
        \b4_nUAi[370] , \b4_nUAi[369] , \b4_nUAi[368] , \b4_nUAi[367] , 
        \b4_nUAi[366] , \b4_nUAi[365] , \b4_nUAi[364] , \b4_nUAi[363] , 
        \b4_nUAi[362] , \b4_nUAi[361] , \b4_nUAi[360] , \b4_nUAi[359] , 
        \b4_nUAi[358] , \b4_nUAi[357] , \b4_nUAi[356] , \b4_nUAi[355] , 
        \b4_nUAi[354] , \b4_nUAi[353] , \b4_nUAi[352] , \b4_nUAi[351] , 
        \b4_nUAi[350] , \b4_nUAi[349] , \b4_nUAi[348] , \b4_nUAi[347] , 
        \b4_nUAi[346] , \b4_nUAi[345] , \b4_nUAi[344] , \b4_nUAi[343] , 
        \b4_nUAi[342] , \b4_nUAi[341] , \b4_nUAi[340] , \b4_nUAi[339] , 
        \b4_nUAi[338] , \b4_nUAi[337] , \b4_nUAi[336] , \b4_nUAi[335] , 
        \b4_nUAi[334] , \b4_nUAi[333] , \b4_nUAi[332] , \b4_nUAi[331] , 
        \b4_nUAi[330] , \b4_nUAi[329] , \b4_nUAi[328] , \b4_nUAi[327] , 
        \b4_nUAi[326] , \b4_nUAi[325] , \b4_nUAi[324] , \b4_nUAi[323] , 
        \b4_nUAi[322] , \b4_nUAi[321] , \b4_nUAi[320] , \b4_nUAi[319] , 
        \b4_nUAi[318] , \b4_nUAi[317] , \b4_nUAi[316] , \b4_nUAi[315] , 
        \b4_nUAi[314] , \b4_nUAi[313] , \b4_nUAi[312] , \b4_nUAi[311] , 
        \b4_nUAi[310] , \b4_nUAi[309] , \b4_nUAi[308] , \b4_nUAi[307] , 
        \b4_nUAi[306] , \b4_nUAi[305] , \b4_nUAi[304] , \b4_nUAi[303] , 
        \b4_nUAi[302] , \b4_nUAi[301] , \b4_nUAi[300] , \b4_nUAi[299] , 
        \b4_nUAi[298] , \b4_nUAi[297] , \b4_nUAi[296] , \b4_nUAi[295] , 
        \b4_nUAi[294] , \b4_nUAi[293] , \b4_nUAi[292] , \b4_nUAi[291] , 
        \b4_nUAi[290] , \b4_nUAi[289] , \b4_nUAi[288] , \b4_nUAi[287] , 
        \b4_nUAi[286] , \b4_nUAi[285] , \b4_nUAi[284] , \b4_nUAi[283] , 
        \b4_nUAi[282] , \b4_nUAi[281] , \b4_nUAi[280] , \b4_nUAi[279] , 
        \b4_nUAi[278] , \b4_nUAi[277] , \b4_nUAi[276] , \b4_nUAi[275] , 
        \b4_nUAi[274] , \b4_nUAi[273] , \b4_nUAi[272] , \b4_nUAi[271] , 
        \b4_nUAi[270] , \b4_nUAi[269] , \b4_nUAi[268] , \b4_nUAi[267] , 
        \b4_nUAi[266] , \b4_nUAi[265] , \b4_nUAi[264] , \b4_nUAi[263] , 
        \b4_nUAi[262] , \b4_nUAi[261] , \b4_nUAi[260] , \b4_nUAi[259] , 
        \b4_nUAi[258] , \b4_nUAi[257] , \b4_nUAi[256] , \b4_nUAi[255] , 
        \b4_nUAi[254] , \b4_nUAi[253] , \b4_nUAi[252] , \b4_nUAi[251] , 
        \b4_nUAi[250] , \b4_nUAi[249] , \b4_nUAi[248] , \b4_nUAi[247] , 
        \b4_nUAi[246] , \b4_nUAi[245] , \b4_nUAi[244] , \b4_nUAi[243] , 
        \b4_nUAi[242] , \b4_nUAi[241] , \b4_nUAi[240] , \b4_nUAi[239] , 
        \b4_nUAi[238] , \b4_nUAi[237] , \b4_nUAi[236] , \b4_nUAi[235] , 
        \b4_nUAi[234] , \b4_nUAi[233] , \b4_nUAi[232] , \b4_nUAi[231] , 
        \b4_nUAi[230] , \b4_nUAi[229] , \b4_nUAi[228] , \b4_nUAi[227] , 
        \b4_nUAi[226] , \b4_nUAi[225] , \b4_nUAi[224] , \b4_nUAi[223] , 
        \b4_nUAi[222] , \b4_nUAi[221] , \b4_nUAi[220] , \b4_nUAi[219] , 
        \b4_nUAi[218] , \b4_nUAi[217] , \b4_nUAi[216] , \b4_nUAi[215] , 
        \b4_nUAi[214] , \b4_nUAi[213] , \b4_nUAi[212] , \b4_nUAi[211] , 
        \b4_nUAi[210] , \b4_nUAi[209] , \b4_nUAi[208] , \b4_nUAi[207] , 
        \b4_nUAi[206] , \b4_nUAi[205] , \b4_nUAi[204] , \b4_nUAi[203] , 
        \b4_nUAi[202] , \b4_nUAi[201] , \b4_nUAi[200] , \b4_nUAi[199] , 
        \b4_nUAi[198] , \b4_nUAi[197] , \b4_nUAi[196] , \b4_nUAi[195] , 
        \b4_nUAi[194] , \b4_nUAi[193] , \b4_nUAi[192] , \b4_nUAi[191] , 
        \b4_nUAi[190] , \b4_nUAi[189] , \b4_nUAi[188] , \b4_nUAi[187] , 
        \b4_nUAi[186] , \b4_nUAi[185] , \b4_nUAi[184] , \b4_nUAi[183] , 
        \b4_nUAi[182] , \b4_nUAi[181] , \b4_nUAi[180] , \b4_nUAi[179] , 
        \b4_nUAi[178] , \b4_nUAi[177] , \b4_nUAi[176] , \b4_nUAi[175] , 
        \b4_nUAi[174] , \b4_nUAi[173] , \b4_nUAi[172] , \b4_nUAi[171] , 
        \b4_nUAi[170] , \b4_nUAi[169] , \b4_nUAi[168] , \b4_nUAi[167] , 
        \b4_nUAi[166] , \b4_nUAi[165] , \b4_nUAi[164] , \b4_nUAi[163] , 
        \b4_nUAi[162] , \b4_nUAi[161] , \b4_nUAi[160] , \b4_nUAi[159] , 
        \b4_nUAi[158] , \b4_nUAi[157] , \b4_nUAi[156] , \b4_nUAi[155] , 
        \b4_nUAi[154] , \b4_nUAi[153] , \b4_nUAi[152] , \b4_nUAi[151] , 
        \b4_nUAi[150] , \b4_nUAi[149] , \b4_nUAi[148] , \b4_nUAi[147] , 
        \b4_nUAi[146] , \b4_nUAi[145] , \b4_nUAi[144] , \b4_nUAi[143] , 
        \b4_nUAi[142] , \b4_nUAi[141] , \b4_nUAi[140] , \b4_nUAi[139] , 
        \b4_nUAi[138] , \b4_nUAi[137] , \b4_nUAi[136] , \b4_nUAi[135] , 
        \b4_nUAi[134] , \b4_nUAi[133] , \b4_nUAi[132] , \b4_nUAi[131] , 
        \b4_nUAi[130] , \b4_nUAi[129] , \b4_nUAi[128] , \b4_nUAi[127] , 
        \b4_nUAi[126] , \b4_nUAi[125] , \b4_nUAi[124] , \b4_nUAi[123] , 
        \b4_nUAi[122] , \b4_nUAi[121] , \b4_nUAi[120] , \b4_nUAi[119] , 
        \b4_nUAi[118] , \b4_nUAi[117] , \b4_nUAi[116] , \b4_nUAi[115] , 
        \b4_nUAi[114] , \b4_nUAi[113] , \b4_nUAi[112] , \b4_nUAi[111] , 
        \b4_nUAi[110] , \b4_nUAi[109] , \b4_nUAi[108] , \b4_nUAi[107] , 
        \b4_nUAi[106] , \b4_nUAi[105] , \b4_nUAi[104] , \b4_nUAi[103] , 
        \b4_nUAi[102] , \b4_nUAi[101] , \b4_nUAi[100] , \b4_nUAi[99] , 
        \b4_nUAi[98] , \b4_nUAi[97] , \b4_nUAi[96] , \b4_nUAi[95] , 
        \b4_nUAi[94] , \b4_nUAi[93] , \b4_nUAi[92] , \b4_nUAi[91] , 
        \b4_nUAi[90] , \b4_nUAi[89] , \b4_nUAi[88] , \b4_nUAi[87] , 
        \b4_nUAi[86] , \b4_nUAi[85] , \b4_nUAi[84] , \b4_nUAi[83] , 
        \b4_nUAi[82] , \b4_nUAi[81] , \b4_nUAi[80] , \b4_nUAi[79] , 
        \b4_nUAi[78] , \b4_nUAi[77] , \b4_nUAi[76] , \b4_nUAi[75] , 
        \b4_nUAi[74] , \b4_nUAi[73] , \b4_nUAi[72] , \b4_nUAi[71] , 
        \b4_nUAi[70] , \b4_nUAi[69] , \b4_nUAi[68] , \b4_nUAi[67] , 
        \b4_nUAi[66] , \b4_nUAi[65] , \b4_nUAi[64] , \b4_nUAi[63] , 
        \b4_nUAi[62] , \b4_nUAi[61] , \b4_nUAi[60] , \b4_nUAi[59] , 
        \b4_nUAi[58] , \b4_nUAi[57] , \b4_nUAi[56] , \b4_nUAi[55] , 
        \b4_nUAi[54] , \b4_nUAi[53] , \b4_nUAi[52] , \b4_nUAi[51] , 
        \b4_nUAi[50] , \b4_nUAi[49] , \b4_nUAi[48] , \b4_nUAi[47] , 
        \b4_nUAi[46] , \b4_nUAi[45] , \b4_nUAi[44] , \b4_nUAi[43] , 
        \b4_nUAi[42] , \b4_nUAi[41] , \b4_nUAi[40] , \b4_nUAi[39] , 
        \b4_nUAi[38] , \b4_nUAi[37] , \b4_nUAi[36] , \b4_nUAi[35] , 
        \b4_nUAi[34] , \b4_nUAi[33] , \b4_nUAi[32] , \b4_nUAi[31] , 
        \b4_nUAi[30] , \b4_nUAi[29] , \b4_nUAi[28] , \b4_nUAi[27] , 
        \b4_nUAi[26] , \b4_nUAi[25] , \b4_nUAi[24] , \b4_nUAi[23] , 
        \b4_nUAi[22] , \b4_nUAi[21] , \b4_nUAi[20] , \b4_nUAi[19] , 
        \b4_nUAi[18] , \b4_nUAi[17] , \b4_nUAi[16] , \b4_nUAi[15] , 
        \b4_nUAi[14] , \b4_nUAi[13] , \b4_nUAi[12] , \b4_nUAi[11] , 
        \b4_nUAi[10] , \b4_nUAi[9] , \b4_nUAi[8] , \b4_nUAi[7] , 
        \b4_nUAi[6] , \b4_nUAi[5] , \b4_nUAi[4] , \b4_nUAi[3] , 
        \b4_nUAi[2] , \b4_nUAi[1] , \b4_nUAi[0] }), .IICE_comm2iice({
        IICE_comm2iice[11], IICE_comm2iice[10]}), .b4_PLyF(b4_PLyF), 
        .b7_PSyi3wy(b7_PSyi3wy), .b8_PSyiBgYG(b8_PSyiBgYG));
    VCC VCC (.Y(VCC_net_1));
    b11_PSyil9s1fkT_x b7_PbTtl9G (.mdiclink_reg({mdiclink_reg[154], 
        mdiclink_reg[153], mdiclink_reg[152], mdiclink_reg[151], 
        mdiclink_reg[150], mdiclink_reg[149], mdiclink_reg[148], 
        mdiclink_reg[147], mdiclink_reg[146], mdiclink_reg[145], 
        mdiclink_reg[144], mdiclink_reg[143], mdiclink_reg[142], 
        mdiclink_reg[141], mdiclink_reg[140], mdiclink_reg[139], 
        mdiclink_reg[138], mdiclink_reg[137], mdiclink_reg[136], 
        mdiclink_reg[135], mdiclink_reg[134], mdiclink_reg[133], 
        mdiclink_reg[132], mdiclink_reg[131], mdiclink_reg[130], 
        mdiclink_reg[129], mdiclink_reg[128], mdiclink_reg[127], 
        mdiclink_reg[126], mdiclink_reg[125], mdiclink_reg[124], 
        mdiclink_reg[123], mdiclink_reg[122], mdiclink_reg[121], 
        mdiclink_reg[120], mdiclink_reg[119], mdiclink_reg[118], 
        mdiclink_reg[117], mdiclink_reg[116], mdiclink_reg[115], 
        mdiclink_reg[114], mdiclink_reg[113], mdiclink_reg[112], 
        mdiclink_reg[111], mdiclink_reg[110], mdiclink_reg[109], 
        mdiclink_reg[108], mdiclink_reg[107], mdiclink_reg[106], 
        mdiclink_reg[105], mdiclink_reg[104], mdiclink_reg[103], 
        mdiclink_reg[102], mdiclink_reg[101], mdiclink_reg[100], 
        mdiclink_reg[99], mdiclink_reg[98], mdiclink_reg[97], 
        mdiclink_reg[96], mdiclink_reg[95], mdiclink_reg[94], 
        mdiclink_reg[93], mdiclink_reg[92], mdiclink_reg[91], 
        mdiclink_reg[90], mdiclink_reg[89], mdiclink_reg[88], 
        mdiclink_reg[87], mdiclink_reg[86], mdiclink_reg[85], 
        mdiclink_reg[84], mdiclink_reg[83], mdiclink_reg[82], 
        mdiclink_reg[81], mdiclink_reg[80], mdiclink_reg[79], 
        mdiclink_reg[78], mdiclink_reg[77], mdiclink_reg[76], 
        mdiclink_reg[75], mdiclink_reg[74], mdiclink_reg[73], 
        mdiclink_reg[72], mdiclink_reg[71], mdiclink_reg[70], 
        mdiclink_reg[69], mdiclink_reg[68], mdiclink_reg[67], 
        mdiclink_reg[66], mdiclink_reg[65], mdiclink_reg[64], 
        mdiclink_reg[63], mdiclink_reg[62], mdiclink_reg[61], 
        mdiclink_reg[60], mdiclink_reg[59], mdiclink_reg[58], 
        mdiclink_reg[57], mdiclink_reg[56], mdiclink_reg[55], 
        mdiclink_reg[54], mdiclink_reg[53], mdiclink_reg[52], 
        mdiclink_reg[51], mdiclink_reg[50], mdiclink_reg[49], 
        mdiclink_reg[48], mdiclink_reg[47], mdiclink_reg[46], 
        mdiclink_reg[45], mdiclink_reg[44], mdiclink_reg[43], 
        mdiclink_reg[42], mdiclink_reg[41], mdiclink_reg[40], 
        mdiclink_reg[39], mdiclink_reg[38], mdiclink_reg[37], 
        mdiclink_reg[36], mdiclink_reg[35], mdiclink_reg[34], 
        mdiclink_reg[33], mdiclink_reg[32], mdiclink_reg[31], 
        mdiclink_reg[30], mdiclink_reg[29], mdiclink_reg[28], 
        mdiclink_reg[27], mdiclink_reg[26], mdiclink_reg[25], 
        mdiclink_reg[24], mdiclink_reg[23], mdiclink_reg[22], 
        mdiclink_reg[21], mdiclink_reg[20], mdiclink_reg[19], 
        mdiclink_reg[18], mdiclink_reg[17], mdiclink_reg[16], 
        mdiclink_reg[15], mdiclink_reg[14], mdiclink_reg[13], 
        mdiclink_reg[12], mdiclink_reg[11], mdiclink_reg[10], 
        mdiclink_reg[9], mdiclink_reg[8], mdiclink_reg[7], 
        mdiclink_reg[6], mdiclink_reg[5], mdiclink_reg[4], 
        mdiclink_reg[3], mdiclink_reg[2], mdiclink_reg[1], 
        mdiclink_reg[0]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[154], 
        b11_OFWNT9L_8tZ[153], b11_OFWNT9L_8tZ[152], 
        b11_OFWNT9L_8tZ[151], b11_OFWNT9L_8tZ[150], 
        b11_OFWNT9L_8tZ[149], b11_OFWNT9L_8tZ[148], 
        b11_OFWNT9L_8tZ[147], b11_OFWNT9L_8tZ[146], 
        b11_OFWNT9L_8tZ[145], b11_OFWNT9L_8tZ[144], 
        b11_OFWNT9L_8tZ[143], b11_OFWNT9L_8tZ[142], 
        b11_OFWNT9L_8tZ[141], b11_OFWNT9L_8tZ[140], 
        b11_OFWNT9L_8tZ[139], b11_OFWNT9L_8tZ[138], 
        b11_OFWNT9L_8tZ[137], b11_OFWNT9L_8tZ[136], 
        b11_OFWNT9L_8tZ[135], b11_OFWNT9L_8tZ[134], 
        b11_OFWNT9L_8tZ[133], b11_OFWNT9L_8tZ[132], 
        b11_OFWNT9L_8tZ[131], b11_OFWNT9L_8tZ[130], 
        b11_OFWNT9L_8tZ[129], b11_OFWNT9L_8tZ[128], 
        b11_OFWNT9L_8tZ[127], b11_OFWNT9L_8tZ[126], 
        b11_OFWNT9L_8tZ[125], b11_OFWNT9L_8tZ[124], 
        b11_OFWNT9L_8tZ[123], b11_OFWNT9L_8tZ[122], 
        b11_OFWNT9L_8tZ[121], b11_OFWNT9L_8tZ[120], 
        b11_OFWNT9L_8tZ[119], b11_OFWNT9L_8tZ[118], 
        b11_OFWNT9L_8tZ[117], b11_OFWNT9L_8tZ[116], 
        b11_OFWNT9L_8tZ[115], b11_OFWNT9L_8tZ[114], 
        b11_OFWNT9L_8tZ[113], b11_OFWNT9L_8tZ[112], 
        b11_OFWNT9L_8tZ[111], b11_OFWNT9L_8tZ[110], 
        b11_OFWNT9L_8tZ[109], b11_OFWNT9L_8tZ[108], 
        b11_OFWNT9L_8tZ[107], b11_OFWNT9L_8tZ[106], 
        b11_OFWNT9L_8tZ[105], b11_OFWNT9L_8tZ[104], 
        b11_OFWNT9L_8tZ[103], b11_OFWNT9L_8tZ[102], 
        b11_OFWNT9L_8tZ[101], b11_OFWNT9L_8tZ[100], 
        b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], b11_OFWNT9L_8tZ[97], 
        b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], b11_OFWNT9L_8tZ[94], 
        b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], b11_OFWNT9L_8tZ[91], 
        b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], b11_OFWNT9L_8tZ[88], 
        b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], b11_OFWNT9L_8tZ[85], 
        b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], b11_OFWNT9L_8tZ[82], 
        b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], b11_OFWNT9L_8tZ[79], 
        b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], b11_OFWNT9L_8tZ[76], 
        b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], b11_OFWNT9L_8tZ[73], 
        b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], b11_OFWNT9L_8tZ[70], 
        b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], b11_OFWNT9L_8tZ[67], 
        b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], b11_OFWNT9L_8tZ[64], 
        b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], b11_OFWNT9L_8tZ[61], 
        b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], b11_OFWNT9L_8tZ[58], 
        b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], b11_OFWNT9L_8tZ[55], 
        b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], b11_OFWNT9L_8tZ[52], 
        b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], b11_OFWNT9L_8tZ[49], 
        b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], b11_OFWNT9L_8tZ[46], 
        b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], b11_OFWNT9L_8tZ[43], 
        b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], b11_OFWNT9L_8tZ[40], 
        b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], b11_OFWNT9L_8tZ[37], 
        b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], b11_OFWNT9L_8tZ[34], 
        b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], b11_OFWNT9L_8tZ[31], 
        b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], b11_OFWNT9L_8tZ[28], 
        b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], b11_OFWNT9L_8tZ[25], 
        b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], b11_OFWNT9L_8tZ[22], 
        b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], b11_OFWNT9L_8tZ[19], 
        b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], b11_OFWNT9L_8tZ[16], 
        b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], b11_OFWNT9L_8tZ[13], 
        b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], b11_OFWNT9L_8tZ[10], 
        b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], b11_OFWNT9L_8tZ[7], 
        b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], b11_OFWNT9L_8tZ[4], 
        b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], b11_OFWNT9L_8tZ[1], 
        b11_OFWNT9L_8tZ[0]}), .b4_nUAi({\b4_nUAi[463] , \b4_nUAi[462] , 
        \b4_nUAi[461] , \b4_nUAi[460] , \b4_nUAi[459] , \b4_nUAi[458] , 
        \b4_nUAi[457] , \b4_nUAi[456] , \b4_nUAi[455] , \b4_nUAi[454] , 
        \b4_nUAi[453] , \b4_nUAi[452] , \b4_nUAi[451] , \b4_nUAi[450] , 
        \b4_nUAi[449] , \b4_nUAi[448] , \b4_nUAi[447] , \b4_nUAi[446] , 
        \b4_nUAi[445] , \b4_nUAi[444] , \b4_nUAi[443] , \b4_nUAi[442] , 
        \b4_nUAi[441] , \b4_nUAi[440] , \b4_nUAi[439] , \b4_nUAi[438] , 
        \b4_nUAi[437] , \b4_nUAi[436] , \b4_nUAi[435] , \b4_nUAi[434] , 
        \b4_nUAi[433] , \b4_nUAi[432] , \b4_nUAi[431] , \b4_nUAi[430] , 
        \b4_nUAi[429] , \b4_nUAi[428] , \b4_nUAi[427] , \b4_nUAi[426] , 
        \b4_nUAi[425] , \b4_nUAi[424] , \b4_nUAi[423] , \b4_nUAi[422] , 
        \b4_nUAi[421] , \b4_nUAi[420] , \b4_nUAi[419] , \b4_nUAi[418] , 
        \b4_nUAi[417] , \b4_nUAi[416] , \b4_nUAi[415] , \b4_nUAi[414] , 
        \b4_nUAi[413] , \b4_nUAi[412] , \b4_nUAi[411] , \b4_nUAi[410] , 
        \b4_nUAi[409] , \b4_nUAi[408] , \b4_nUAi[407] , \b4_nUAi[406] , 
        \b4_nUAi[405] , \b4_nUAi[404] , \b4_nUAi[403] , \b4_nUAi[402] , 
        \b4_nUAi[401] , \b4_nUAi[400] , \b4_nUAi[399] , \b4_nUAi[398] , 
        \b4_nUAi[397] , \b4_nUAi[396] , \b4_nUAi[395] , \b4_nUAi[394] , 
        \b4_nUAi[393] , \b4_nUAi[392] , \b4_nUAi[391] , \b4_nUAi[390] , 
        \b4_nUAi[389] , \b4_nUAi[388] , \b4_nUAi[387] , \b4_nUAi[386] , 
        \b4_nUAi[385] , \b4_nUAi[384] , \b4_nUAi[383] , \b4_nUAi[382] , 
        \b4_nUAi[381] , \b4_nUAi[380] , \b4_nUAi[379] , \b4_nUAi[378] , 
        \b4_nUAi[377] , \b4_nUAi[376] , \b4_nUAi[375] , \b4_nUAi[374] , 
        \b4_nUAi[373] , \b4_nUAi[372] , \b4_nUAi[371] , \b4_nUAi[370] , 
        \b4_nUAi[369] , \b4_nUAi[368] , \b4_nUAi[367] , \b4_nUAi[366] , 
        \b4_nUAi[365] , \b4_nUAi[364] , \b4_nUAi[363] , \b4_nUAi[362] , 
        \b4_nUAi[361] , \b4_nUAi[360] , \b4_nUAi[359] , \b4_nUAi[358] , 
        \b4_nUAi[357] , \b4_nUAi[356] , \b4_nUAi[355] , \b4_nUAi[354] , 
        \b4_nUAi[353] , \b4_nUAi[352] , \b4_nUAi[351] , \b4_nUAi[350] , 
        \b4_nUAi[349] , \b4_nUAi[348] , \b4_nUAi[347] , \b4_nUAi[346] , 
        \b4_nUAi[345] , \b4_nUAi[344] , \b4_nUAi[343] , \b4_nUAi[342] , 
        \b4_nUAi[341] , \b4_nUAi[340] , \b4_nUAi[339] , \b4_nUAi[338] , 
        \b4_nUAi[337] , \b4_nUAi[336] , \b4_nUAi[335] , \b4_nUAi[334] , 
        \b4_nUAi[333] , \b4_nUAi[332] , \b4_nUAi[331] , \b4_nUAi[330] , 
        \b4_nUAi[329] , \b4_nUAi[328] , \b4_nUAi[327] , \b4_nUAi[326] , 
        \b4_nUAi[325] , \b4_nUAi[324] , \b4_nUAi[323] , \b4_nUAi[322] , 
        \b4_nUAi[321] , \b4_nUAi[320] , \b4_nUAi[319] , \b4_nUAi[318] , 
        \b4_nUAi[317] , \b4_nUAi[316] , \b4_nUAi[315] , \b4_nUAi[314] , 
        \b4_nUAi[313] , \b4_nUAi[312] , \b4_nUAi[311] , \b4_nUAi[310] , 
        \b4_nUAi[309] , \b4_nUAi[308] , \b4_nUAi[307] , \b4_nUAi[306] , 
        \b4_nUAi[305] , \b4_nUAi[304] , \b4_nUAi[303] , \b4_nUAi[302] , 
        \b4_nUAi[301] , \b4_nUAi[300] , \b4_nUAi[299] , \b4_nUAi[298] , 
        \b4_nUAi[297] , \b4_nUAi[296] , \b4_nUAi[295] , \b4_nUAi[294] , 
        \b4_nUAi[293] , \b4_nUAi[292] , \b4_nUAi[291] , \b4_nUAi[290] , 
        \b4_nUAi[289] , \b4_nUAi[288] , \b4_nUAi[287] , \b4_nUAi[286] , 
        \b4_nUAi[285] , \b4_nUAi[284] , \b4_nUAi[283] , \b4_nUAi[282] , 
        \b4_nUAi[281] , \b4_nUAi[280] , \b4_nUAi[279] , \b4_nUAi[278] , 
        \b4_nUAi[277] , \b4_nUAi[276] , \b4_nUAi[275] , \b4_nUAi[274] , 
        \b4_nUAi[273] , \b4_nUAi[272] , \b4_nUAi[271] , \b4_nUAi[270] , 
        \b4_nUAi[269] , \b4_nUAi[268] , \b4_nUAi[267] , \b4_nUAi[266] , 
        \b4_nUAi[265] , \b4_nUAi[264] , \b4_nUAi[263] , \b4_nUAi[262] , 
        \b4_nUAi[261] , \b4_nUAi[260] , \b4_nUAi[259] , \b4_nUAi[258] , 
        \b4_nUAi[257] , \b4_nUAi[256] , \b4_nUAi[255] , \b4_nUAi[254] , 
        \b4_nUAi[253] , \b4_nUAi[252] , \b4_nUAi[251] , \b4_nUAi[250] , 
        \b4_nUAi[249] , \b4_nUAi[248] , \b4_nUAi[247] , \b4_nUAi[246] , 
        \b4_nUAi[245] , \b4_nUAi[244] , \b4_nUAi[243] , \b4_nUAi[242] , 
        \b4_nUAi[241] , \b4_nUAi[240] , \b4_nUAi[239] , \b4_nUAi[238] , 
        \b4_nUAi[237] , \b4_nUAi[236] , \b4_nUAi[235] , \b4_nUAi[234] , 
        \b4_nUAi[233] , \b4_nUAi[232] , \b4_nUAi[231] , \b4_nUAi[230] , 
        \b4_nUAi[229] , \b4_nUAi[228] , \b4_nUAi[227] , \b4_nUAi[226] , 
        \b4_nUAi[225] , \b4_nUAi[224] , \b4_nUAi[223] , \b4_nUAi[222] , 
        \b4_nUAi[221] , \b4_nUAi[220] , \b4_nUAi[219] , \b4_nUAi[218] , 
        \b4_nUAi[217] , \b4_nUAi[216] , \b4_nUAi[215] , \b4_nUAi[214] , 
        \b4_nUAi[213] , \b4_nUAi[212] , \b4_nUAi[211] , \b4_nUAi[210] , 
        \b4_nUAi[209] , \b4_nUAi[208] , \b4_nUAi[207] , \b4_nUAi[206] , 
        \b4_nUAi[205] , \b4_nUAi[204] , \b4_nUAi[203] , \b4_nUAi[202] , 
        \b4_nUAi[201] , \b4_nUAi[200] , \b4_nUAi[199] , \b4_nUAi[198] , 
        \b4_nUAi[197] , \b4_nUAi[196] , \b4_nUAi[195] , \b4_nUAi[194] , 
        \b4_nUAi[193] , \b4_nUAi[192] , \b4_nUAi[191] , \b4_nUAi[190] , 
        \b4_nUAi[189] , \b4_nUAi[188] , \b4_nUAi[187] , \b4_nUAi[186] , 
        \b4_nUAi[185] , \b4_nUAi[184] , \b4_nUAi[183] , \b4_nUAi[182] , 
        \b4_nUAi[181] , \b4_nUAi[180] , \b4_nUAi[179] , \b4_nUAi[178] , 
        \b4_nUAi[177] , \b4_nUAi[176] , \b4_nUAi[175] , \b4_nUAi[174] , 
        \b4_nUAi[173] , \b4_nUAi[172] , \b4_nUAi[171] , \b4_nUAi[170] , 
        \b4_nUAi[169] , \b4_nUAi[168] , \b4_nUAi[167] , \b4_nUAi[166] , 
        \b4_nUAi[165] , \b4_nUAi[164] , \b4_nUAi[163] , \b4_nUAi[162] , 
        \b4_nUAi[161] , \b4_nUAi[160] , \b4_nUAi[159] , \b4_nUAi[158] , 
        \b4_nUAi[157] , \b4_nUAi[156] , \b4_nUAi[155] , \b4_nUAi[154] , 
        \b4_nUAi[153] , \b4_nUAi[152] , \b4_nUAi[151] , \b4_nUAi[150] , 
        \b4_nUAi[149] , \b4_nUAi[148] , \b4_nUAi[147] , \b4_nUAi[146] , 
        \b4_nUAi[145] , \b4_nUAi[144] , \b4_nUAi[143] , \b4_nUAi[142] , 
        \b4_nUAi[141] , \b4_nUAi[140] , \b4_nUAi[139] , \b4_nUAi[138] , 
        \b4_nUAi[137] , \b4_nUAi[136] , \b4_nUAi[135] , \b4_nUAi[134] , 
        \b4_nUAi[133] , \b4_nUAi[132] , \b4_nUAi[131] , \b4_nUAi[130] , 
        \b4_nUAi[129] , \b4_nUAi[128] , \b4_nUAi[127] , \b4_nUAi[126] , 
        \b4_nUAi[125] , \b4_nUAi[124] , \b4_nUAi[123] , \b4_nUAi[122] , 
        \b4_nUAi[121] , \b4_nUAi[120] , \b4_nUAi[119] , \b4_nUAi[118] , 
        \b4_nUAi[117] , \b4_nUAi[116] , \b4_nUAi[115] , \b4_nUAi[114] , 
        \b4_nUAi[113] , \b4_nUAi[112] , \b4_nUAi[111] , \b4_nUAi[110] , 
        \b4_nUAi[109] , \b4_nUAi[108] , \b4_nUAi[107] , \b4_nUAi[106] , 
        \b4_nUAi[105] , \b4_nUAi[104] , \b4_nUAi[103] , \b4_nUAi[102] , 
        \b4_nUAi[101] , \b4_nUAi[100] , \b4_nUAi[99] , \b4_nUAi[98] , 
        \b4_nUAi[97] , \b4_nUAi[96] , \b4_nUAi[95] , \b4_nUAi[94] , 
        \b4_nUAi[93] , \b4_nUAi[92] , \b4_nUAi[91] , \b4_nUAi[90] , 
        \b4_nUAi[89] , \b4_nUAi[88] , \b4_nUAi[87] , \b4_nUAi[86] , 
        \b4_nUAi[85] , \b4_nUAi[84] , \b4_nUAi[83] , \b4_nUAi[82] , 
        \b4_nUAi[81] , \b4_nUAi[80] , \b4_nUAi[79] , \b4_nUAi[78] , 
        \b4_nUAi[77] , \b4_nUAi[76] , \b4_nUAi[75] , \b4_nUAi[74] , 
        \b4_nUAi[73] , \b4_nUAi[72] , \b4_nUAi[71] , \b4_nUAi[70] , 
        \b4_nUAi[69] , \b4_nUAi[68] , \b4_nUAi[67] , \b4_nUAi[66] , 
        \b4_nUAi[65] , \b4_nUAi[64] , \b4_nUAi[63] , \b4_nUAi[62] , 
        \b4_nUAi[61] , \b4_nUAi[60] , \b4_nUAi[59] , \b4_nUAi[58] , 
        \b4_nUAi[57] , \b4_nUAi[56] , \b4_nUAi[55] , \b4_nUAi[54] , 
        \b4_nUAi[53] , \b4_nUAi[52] , \b4_nUAi[51] , \b4_nUAi[50] , 
        \b4_nUAi[49] , \b4_nUAi[48] , \b4_nUAi[47] , \b4_nUAi[46] , 
        \b4_nUAi[45] , \b4_nUAi[44] , \b4_nUAi[43] , \b4_nUAi[42] , 
        \b4_nUAi[41] , \b4_nUAi[40] , \b4_nUAi[39] , \b4_nUAi[38] , 
        \b4_nUAi[37] , \b4_nUAi[36] , \b4_nUAi[35] , \b4_nUAi[34] , 
        \b4_nUAi[33] , \b4_nUAi[32] , \b4_nUAi[31] , \b4_nUAi[30] , 
        \b4_nUAi[29] , \b4_nUAi[28] , \b4_nUAi[27] , \b4_nUAi[26] , 
        \b4_nUAi[25] , \b4_nUAi[24] , \b4_nUAi[23] , \b4_nUAi[22] , 
        \b4_nUAi[21] , \b4_nUAi[20] , \b4_nUAi[19] , \b4_nUAi[18] , 
        \b4_nUAi[17] , \b4_nUAi[16] , \b4_nUAi[15] , \b4_nUAi[14] , 
        \b4_nUAi[13] , \b4_nUAi[12] , \b4_nUAi[11] , \b4_nUAi[10] , 
        \b4_nUAi[9] , \b4_nUAi[8] , \b4_nUAi[7] , \b4_nUAi[6] , 
        \b4_nUAi[5] , \b4_nUAi[4] , \b4_nUAi[3] , \b4_nUAi[2] , 
        \b4_nUAi[1] , \b4_nUAi[0] }), .b11_uUT0JC4gFrY({
        \b11_uUT0JC4gFrY[1] }), .b7_PSyi3wy(b7_PSyi3wy), .BW_clk_c(
        BW_clk_c));
    GND GND (.Y(GND_net_1));
    SLE b7_PSyil9s (.D(\b11_uUT0JC4gFrY[1] ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b11_PSyil9s_FMZ));
    
endmodule


module b8_nR_ymqrG_10s_5s_0_0s_0s_1_510_x_0(
       b6_nfs_IF_i_0,
       b6_nUT_IF,
       b6_nfs_IF,
       IICE_comm2iice_3,
       IICE_comm2iice_0,
       IICE_comm2iice_2,
       b4_PLyF,
       b13_nUTQBgfDb_Z4D,
       b12_nUTQBgfDb_bd,
       b16_nYhI39swMeEd_A78,
       b15_nYhI39swMeEd_Mg,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_qH,
       b11_vABZ3qsY_XH
    );
output [1:1] b6_nfs_IF_i_0;
output [9:0] b6_nUT_IF;
output [4:0] b6_nfs_IF;
input  IICE_comm2iice_3;
input  IICE_comm2iice_0;
input  IICE_comm2iice_2;
input  b4_PLyF;
output b13_nUTQBgfDb_Z4D;
input  b12_nUTQBgfDb_bd;
output b16_nYhI39swMeEd_A78;
input  b15_nYhI39swMeEd_Mg;
output b12_vABZ3qsY_Lyh;
output b11_vABZ3qsY_qH;
input  b11_vABZ3qsY_XH;

    wire \b10_nUT_M9kYfr[2]_net_1 , VCC_net_1, 
        \b10_nUT_M9kYfr[3]_net_1 , b10_nUT_M9kYfr4_net_1, GND_net_1, 
        \b10_nUT_M9kYfr[4]_net_1 , \b10_nUT_M9kYfr[5]_net_1 , 
        \b10_nUT_M9kYfr[6]_net_1 , \b10_nUT_M9kYfr[7]_net_1 , 
        \b10_nUT_M9kYfr[8]_net_1 , \b10_nUT_M9kYfr[9]_net_1 , 
        \b10_nfs_M9kYfr[1]_net_1 , b10_nfs_M9kYfr4_net_1, 
        \b10_nfs_M9kYfr[2]_net_1 , \b10_nfs_M9kYfr[3]_net_1 , 
        \b10_nfs_M9kYfr[4]_net_1 , \b10_nUT_M9kYfr[1]_net_1 , 
        b15_vABZ3qsY_ub3Rme3_net_1, b8_vABZ3qsY_RNO;
    
    SLE \genblk1.b3_nfs[4]  (.D(\b10_nfs_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[4]));
    SLE \b10_nUT_M9kYfr[6]  (.D(\b10_nUT_M9kYfr[7]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[6]_net_1 ));
    SLE \genblk2.b3_nUT[9]  (.D(\b10_nUT_M9kYfr[9]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[9]));
    CFG1 #( .INIT(2'h1) )  \genblk1.b3_nfs_RNI8HD5[1]  (.A(
        b6_nfs_IF[1]), .Y(b6_nfs_IF_i_0[1]));
    SLE \genblk2.b3_nUT[6]  (.D(\b10_nUT_M9kYfr[6]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[6]));
    SLE \b10_nUT_M9kYfr[9]  (.D(b4_PLyF), .CLK(IICE_comm2iice_3), .EN(
        b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b10_nUT_M9kYfr[9]_net_1 ));
    CFG2 #( .INIT(4'h8) )  b10_nfs_M9kYfr4 (.A(b12_nUTQBgfDb_bd), .B(
        IICE_comm2iice_2), .Y(b10_nfs_M9kYfr4_net_1));
    SLE \genblk2.b3_nUT[3]  (.D(\b10_nUT_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[3]));
    SLE \b10_nfs_M9kYfr[2]  (.D(\b10_nfs_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nfs_M9kYfr[2]_net_1 ));
    SLE \genblk2.b3_nUT[2]  (.D(\b10_nUT_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[2]));
    SLE \b10_nUT_M9kYfr[3]  (.D(\b10_nUT_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[3]_net_1 ));
    SLE b15_vABZ3qsY_ub3Rme (.D(b4_PLyF), .CLK(IICE_comm2iice_3), .EN(
        b15_vABZ3qsY_ub3Rme3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b12_vABZ3qsY_Lyh));
    VCC VCC (.Y(VCC_net_1));
    SLE \b10_nfs_M9kYfr[3]  (.D(\b10_nfs_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nfs_M9kYfr[3]_net_1 ));
    SLE \genblk1.b3_nfs[3]  (.D(\b10_nfs_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[3]));
    SLE \genblk2.b3_nUT[7]  (.D(\b10_nUT_M9kYfr[7]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[7]));
    SLE \genblk1.b3_nfs[1]  (.D(\b10_nfs_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[1]));
    SLE \b10_nfs_M9kYfr[1]  (.D(\b10_nfs_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nfs_M9kYfr[1]_net_1 ));
    SLE \b10_nUT_M9kYfr[4]  (.D(\b10_nUT_M9kYfr[5]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[4]_net_1 ));
    SLE \genblk2.b3_nUT[0]  (.D(b16_nYhI39swMeEd_A78), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[0]));
    SLE \b10_nUT_M9kYfr[1]  (.D(\b10_nUT_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[1]_net_1 ));
    SLE \b10_nUT_M9kYfr[0]  (.D(\b10_nUT_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b16_nYhI39swMeEd_A78));
    GND GND (.Y(GND_net_1));
    SLE \genblk2.b3_nUT[8]  (.D(\b10_nUT_M9kYfr[8]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[8]));
    SLE \b10_nfs_M9kYfr[4]  (.D(b4_PLyF), .CLK(IICE_comm2iice_3), .EN(
        b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b10_nfs_M9kYfr[4]_net_1 ));
    SLE \genblk2.b3_nUT[4]  (.D(\b10_nUT_M9kYfr[4]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[4]));
    SLE \b10_nfs_M9kYfr[0]  (.D(\b10_nfs_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nfs_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b13_nUTQBgfDb_Z4D));
    SLE \b10_nUT_M9kYfr[7]  (.D(\b10_nUT_M9kYfr[8]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  b10_nUT_M9kYfr4 (.A(b15_nYhI39swMeEd_Mg), 
        .B(IICE_comm2iice_2), .Y(b10_nUT_M9kYfr4_net_1));
    SLE \b10_nUT_M9kYfr[8]  (.D(\b10_nUT_M9kYfr[9]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[8]_net_1 ));
    SLE \genblk1.b3_nfs[2]  (.D(\b10_nfs_M9kYfr[2]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[2]));
    SLE \genblk1.b3_nfs[0]  (.D(b13_nUTQBgfDb_Z4D), .CLK(
        IICE_comm2iice_0), .EN(b12_nUTQBgfDb_bd), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nfs_IF[0]));
    SLE \genblk3.b8_vABZ3qsY  (.D(b12_vABZ3qsY_Lyh), .CLK(
        IICE_comm2iice_0), .EN(b8_vABZ3qsY_RNO), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b11_vABZ3qsY_qH));
    SLE \b10_nUT_M9kYfr[5]  (.D(\b10_nUT_M9kYfr[6]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[5]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \genblk3.b8_vABZ3qsY_RNO  (.A(
        b11_vABZ3qsY_XH), .B(b6_nfs_IF[1]), .Y(b8_vABZ3qsY_RNO));
    SLE \genblk2.b3_nUT[5]  (.D(\b10_nUT_M9kYfr[5]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[5]));
    CFG2 #( .INIT(4'h8) )  b15_vABZ3qsY_ub3Rme3 (.A(b11_vABZ3qsY_XH), 
        .B(IICE_comm2iice_2), .Y(b15_vABZ3qsY_ub3Rme3_net_1));
    SLE \b10_nUT_M9kYfr[2]  (.D(\b10_nUT_M9kYfr[3]_net_1 ), .CLK(
        IICE_comm2iice_3), .EN(b10_nUT_M9kYfr4_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b10_nUT_M9kYfr[2]_net_1 ));
    SLE \genblk2.b3_nUT[1]  (.D(\b10_nUT_M9kYfr[1]_net_1 ), .CLK(
        IICE_comm2iice_0), .EN(b15_nYhI39swMeEd_Mg), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b6_nUT_IF[1]));
    
endmodule


module clock2_en_reg_en_5s_x_0(
       IICE_comm2iice,
       b6_nfs_IF_i_0,
       status_b2sclk,
       b6_nfs_IF,
       b6_Ocm0rW,
       b13_nAzGfFM_sLsv3_3,
       b13_nAzGfFM_sLsv3_0,
       b13_nAzGfFM_sLsv3_2,
       BW_clk_c,
       N_38,
       N_78
    );
input  [11:11] IICE_comm2iice;
input  [1:1] b6_nfs_IF_i_0;
output [3:0] status_b2sclk;
input  [1:1] b6_nfs_IF;
input  [2:2] b6_Ocm0rW;
input  b13_nAzGfFM_sLsv3_3;
input  b13_nAzGfFM_sLsv3_0;
input  b13_nAzGfFM_sLsv3_2;
input  BW_clk_c;
input  N_38;
input  N_78;

    wire src_ack_net_1, src_ack_i_0, VCC_net_1, \int_data[0]_net_1 , 
        dout4_0_a2_RNIKLH5_net_1, GND_net_1, \int_data[1]_net_1 , 
        \int_data[2]_net_1 , \int_data[3]_net_1 , dout4, N_61_i_0, 
        in_en_RNICUKI_net_1, N_19_i_0, in_en_net_1, src_req_net_1, 
        src_req_RNO_0_net_1, in_enc_1_i, N_70_i_0, in_enc_net_1, 
        dst_req_d_net_1, dst_req_d_0, dst_req_net_1, dst_req_0;
    
    SLE \dout[1]  (.D(\int_data[1]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[1]));
    CFG2 #( .INIT(4'h4) )  dst_req_r (.A(b6_nfs_IF[1]), .B(
        src_req_net_1), .Y(dst_req_0));
    CFG2 #( .INIT(4'hE) )  src_req_RNO_0 (.A(in_enc_1_i), .B(
        b6_nfs_IF[1]), .Y(src_req_RNO_0_net_1));
    CFG3 #( .INIT(8'hAB) )  \int_data_RNO[1]  (.A(b13_nAzGfFM_sLsv3_2), 
        .B(N_78), .C(N_38), .Y(N_19_i_0));
    SLE \dout[3]  (.D(\int_data[3]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[3]));
    SLE \int_data[1]  (.D(N_19_i_0), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[1]_net_1 ));
    SLE \dout[2]  (.D(\int_data[2]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[2]));
    GND GND (.Y(GND_net_1));
    SLE in_en (.D(in_enc_net_1), .CLK(BW_clk_c), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(b6_nfs_IF_i_0[1]), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(in_en_net_1));
    CFG2 #( .INIT(4'hE) )  src_ack_RNO (.A(dst_req_net_1), .B(
        dst_req_d_net_1), .Y(N_70_i_0));
    SLE src_ack (.D(N_70_i_0), .CLK(BW_clk_c), .EN(VCC_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(b6_nfs_IF_i_0[1]), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(src_ack_net_1));
    SLE \int_data[0]  (.D(N_61_i_0), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[0]_net_1 ));
    SLE \int_data[2]  (.D(b6_Ocm0rW[2]), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[2]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \int_data_RNO[0]  (.A(N_38), .B(
        b13_nAzGfFM_sLsv3_0), .Y(N_61_i_0));
    SLE \dout[0]  (.D(\int_data[0]_net_1 ), .CLK(IICE_comm2iice[11]), 
        .EN(dout4_0_a2_RNIKLH5_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        status_b2sclk[0]));
    CFG2 #( .INIT(4'hE) )  src_req_RNO_1 (.A(in_en_net_1), .B(
        src_ack_net_1), .Y(in_enc_1_i));
    CFG3 #( .INIT(8'h01) )  in_enc (.A(src_req_net_1), .B(
        src_ack_net_1), .C(in_en_net_1), .Y(in_enc_net_1));
    SLE dst_req (.D(dst_req_0), .CLK(IICE_comm2iice[11]), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dst_req_net_1));
    CFG1 #( .INIT(2'h1) )  src_req_RNO (.A(src_ack_net_1), .Y(
        src_ack_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hE) )  in_en_RNICUKI (.A(b6_nfs_IF[1]), .B(
        in_en_net_1), .Y(in_en_RNICUKI_net_1));
    CFG2 #( .INIT(4'h2) )  dout4_0_a2 (.A(dst_req_net_1), .B(
        dst_req_d_net_1), .Y(dout4));
    SLE \int_data[3]  (.D(b13_nAzGfFM_sLsv3_3), .CLK(BW_clk_c), .EN(
        in_en_RNICUKI_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \int_data[3]_net_1 ));
    CFG2 #( .INIT(4'hE) )  dout4_0_a2_RNIKLH5 (.A(b6_nfs_IF[1]), .B(
        dout4), .Y(dout4_0_a2_RNIKLH5_net_1));
    SLE src_req (.D(src_ack_i_0), .CLK(BW_clk_c), .EN(
        src_req_RNO_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b6_nfs_IF_i_0[1]), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        src_req_net_1));
    SLE dst_req_d (.D(dst_req_d_0), .CLK(IICE_comm2iice[11]), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(dst_req_d_net_1));
    CFG2 #( .INIT(4'h4) )  dst_req_d_r (.A(b6_nfs_IF[1]), .B(
        dst_req_net_1), .Y(dst_req_d_0));
    
endmodule


module b7_OCByLXC_Z1_x_0(
       IICE_comm2iice,
       b13_nAzGfFM_sLsv3_0,
       b8_SoWGfWYY,
       b8_SoWGfWYY_i,
       BW_clk_c,
       b12_uRrc2XfY_Lyh,
       N_44,
       b11_PSyil9s_FMZ,
       b4_PLyF,
       b11_uRrc2XfY_XH,
       b13_nUTQBgfDb_Z4D,
       b12_nUTQBgfDb_bd,
       b16_nYhI39swMeEd_A78,
       b15_nYhI39swMeEd_Mg,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_XH
    );
input  [11:8] IICE_comm2iice;
output b13_nAzGfFM_sLsv3_0;
output b8_SoWGfWYY;
output b8_SoWGfWYY_i;
input  BW_clk_c;
output b12_uRrc2XfY_Lyh;
output N_44;
input  b11_PSyil9s_FMZ;
input  b4_PLyF;
input  b11_uRrc2XfY_XH;
output b13_nUTQBgfDb_Z4D;
input  b12_nUTQBgfDb_bd;
output b16_nYhI39swMeEd_A78;
input  b15_nYhI39swMeEd_Mg;
output b12_vABZ3qsY_Lyh;
input  b11_vABZ3qsY_XH;

    wire \b13_nAzGfFM_sLsv3_i[0]_net_1 , \b13_nAzGfFM_sLsv3_i_i_0[0] , 
        \b3_nfs[0]_net_1 , VCC_net_1, \b6_nfs_IF[0] , GND_net_1, 
        \b3_nfs[1]_net_1 , \b6_nfs_IF[1] , \b3_nfs[2]_net_1 , 
        \b6_nfs_IF[2] , \b3_nfs[3]_net_1 , \b6_nfs_IF[3] , 
        \b3_nfs[4]_net_1 , \b6_nfs_IF[4] , 
        \b12_uRrc2XfY_rbN[19]_net_1 , \b12_uRrc2XfY_rbN_5[19]_net_1 , 
        un1_b12_uRrc2XfY_rbN10_i_0, \b12_uRrc2XfY_rbN[20]_net_1 , 
        \b12_uRrc2XfY_rbN_5[20]_net_1 , \b12_uRrc2XfY_rbN[21]_net_1 , 
        \b12_uRrc2XfY_rbN_5[21]_net_1 , \b12_uRrc2XfY_rbN[22]_net_1 , 
        \b12_uRrc2XfY_rbN_5[22]_net_1 , \b12_uRrc2XfY_rbN[23]_net_1 , 
        \b12_uRrc2XfY_rbN_5[23]_net_1 , \b12_uRrc2XfY_rbN[24]_net_1 , 
        \b12_uRrc2XfY_rbN_5[24]_net_1 , \b12_uRrc2XfY_rbN[25]_net_1 , 
        \b12_uRrc2XfY_rbN_5[25]_net_1 , \b12_uRrc2XfY_rbN[4]_net_1 , 
        \b12_uRrc2XfY_rbN_5[4]_net_1 , \b12_uRrc2XfY_rbN[5]_net_1 , 
        \b12_uRrc2XfY_rbN_5[5]_net_1 , \b12_uRrc2XfY_rbN[6]_net_1 , 
        \b12_uRrc2XfY_rbN_5[6]_net_1 , \b12_uRrc2XfY_rbN[7]_net_1 , 
        \b12_uRrc2XfY_rbN_5[7]_net_1 , \b12_uRrc2XfY_rbN[8]_net_1 , 
        \b12_uRrc2XfY_rbN_5[8]_net_1 , \b12_uRrc2XfY_rbN[9]_net_1 , 
        \b12_uRrc2XfY_rbN_5[9]_net_1 , \b12_uRrc2XfY_rbN[10]_net_1 , 
        \b12_uRrc2XfY_rbN_5[10]_net_1 , \b12_uRrc2XfY_rbN[11]_net_1 , 
        \b12_uRrc2XfY_rbN_5[11]_net_1 , \b12_uRrc2XfY_rbN[12]_net_1 , 
        \b12_uRrc2XfY_rbN_5[12]_net_1 , \b12_uRrc2XfY_rbN[13]_net_1 , 
        \b12_uRrc2XfY_rbN_5[13]_net_1 , \b12_uRrc2XfY_rbN[14]_net_1 , 
        \b12_uRrc2XfY_rbN_5[14]_net_1 , \b12_uRrc2XfY_rbN[15]_net_1 , 
        \b12_uRrc2XfY_rbN_5[15]_net_1 , \b12_uRrc2XfY_rbN[16]_net_1 , 
        \b12_uRrc2XfY_rbN_5[16]_net_1 , \b12_uRrc2XfY_rbN[17]_net_1 , 
        \b12_uRrc2XfY_rbN_5[17]_net_1 , \b12_uRrc2XfY_rbN[18]_net_1 , 
        \b12_uRrc2XfY_rbN_5[18]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[15]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[15]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[16]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[16]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[17]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[17]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[18]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[18]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[19]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[19]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[20]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[20]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[21]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[21]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[22]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[22]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[23]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[23]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[24]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[24]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[25]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[25]_net_1 , \b12_uRrc2XfY_rbN_5[0]_net_1 , 
        \b12_uRrc2XfY_rbN[1]_net_1 , \b12_uRrc2XfY_rbN_5[1]_net_1 , 
        \b12_uRrc2XfY_rbN[2]_net_1 , \b12_uRrc2XfY_rbN_5[2]_net_1 , 
        \b12_uRrc2XfY_rbN[3]_net_1 , \b12_uRrc2XfY_rbN_5[3]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[0]_net_1 , \b15_uRrc2XfY_rbN_gr[0]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[1]_net_1 , \b15_uRrc2XfY_rbN_gr[1]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[2]_net_1 , \b15_uRrc2XfY_rbN_gr[2]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[3]_net_1 , \b15_uRrc2XfY_rbN_gr[3]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[5]_net_1 , \b15_uRrc2XfY_rbN_gr[5]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[6]_net_1 , \b15_uRrc2XfY_rbN_gr[6]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[7]_net_1 , \b15_uRrc2XfY_rbN_gr[7]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[8]_net_1 , \b15_uRrc2XfY_rbN_gr[8]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[9]_net_1 , \b15_uRrc2XfY_rbN_gr[9]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[10]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[10]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[11]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[11]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[12]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[12]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[13]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[13]_net_1 , 
        \b15_uRrc2XfY_rbN_gs[14]_net_1 , 
        \b15_uRrc2XfY_rbN_gr[14]_net_1 , N_103_i_0, N_104_i_0, 
        \b13_nAzGfFM_sLsv3[5]_net_1 , b11_vABZ3qsY_qH, 
        \b7_nYhI39s[0]_net_1 , \b7_nYhI39s[1]_net_1 , 
        \b7_nYhI39s[2]_net_1 , \b7_nYhI39s[3]_net_1 , 
        \b7_nYhI39s[4]_net_1 , \b7_nYhI39s[5]_net_1 , 
        \b7_nYhI39s[6]_net_1 , \b7_nYhI39s[7]_net_1 , 
        \b7_nYhI39s[8]_net_1 , \b7_nYhI39s[9]_net_1 , 
        \status_b2sclk[0] , \status_b2sclk[1] , \status_b2sclk[2] , 
        \status_b2sclk[3] , \b13_nAzGfFM_sLsv3[2]_net_1 , 
        \b6_nfs_IF_i_0[1] , N_94_i_0, N_16, 
        \b13_nAzGfFM_sLsv3[3]_net_1 , N_90_i_0, 
        \b13_nAzGfFM_sLsv3[4]_net_1 , N_26_i_0, N_28_i_0, 
        b10_nYhI3_umjB_net_1, b10_nYhI3_umjB_3, 
        un1_b13_nAzGfFM_sLsv3_1_i_0, b8_vABZ3qsY_net_1, 
        \b3_nUT[8]_net_1 , \b6_nUT_IF[8] , \b3_nUT[9]_net_1 , 
        \b6_nUT_IF[9] , \b3_nUT[0]_net_1 , \b6_nUT_IF[0] , 
        \b3_nUT[1]_net_1 , \b6_nUT_IF[1] , \b3_nUT[2]_net_1 , 
        \b6_nUT_IF[2] , \b3_nUT[3]_net_1 , \b6_nUT_IF[3] , 
        \b3_nUT[4]_net_1 , \b6_nUT_IF[4] , \b3_nUT[5]_net_1 , 
        \b6_nUT_IF[5] , \b3_nUT[6]_net_1 , \b6_nUT_IF[6] , 
        \b3_nUT[7]_net_1 , \b6_nUT_IF[7] , \b7_nYhI39s_s[0] , N_23_i_0, 
        \b7_nYhI39s_s[1] , \b7_nYhI39s_s[2] , \b7_nYhI39s_s[3] , 
        \b7_nYhI39s_s[4] , \b7_nYhI39s_s[5] , \b7_nYhI39s_s[6] , 
        \b7_nYhI39s_s[7] , \b7_nYhI39s_s[8] , \b7_nYhI39s_s[9] , 
        b7_nYhI39s_cry_cy, \b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] , N_38, 
        \b7_nYhI39s_cry[0] , \b7_nYhI39s_5[0]_net_1 , 
        \b7_nYhI39s_cry[1] , \b7_nYhI39s_5[1]_net_1 , 
        \b7_nYhI39s_cry[2] , \b7_nYhI39s_5[2]_net_1 , 
        \b7_nYhI39s_cry[3] , \b7_nYhI39s_5[3]_net_1 , 
        \b7_nYhI39s_cry[4] , \b7_nYhI39s_5[4]_net_1 , 
        \b7_nYhI39s_cry[5] , \b7_nYhI39s_5[5]_net_1 , 
        \b7_nYhI39s_cry[6] , \b7_nYhI39s_5[6]_net_1 , 
        \b7_nYhI39s_cry[7] , \b7_nYhI39s_5[7]_net_1 , 
        \b7_nYhI39s_5[9]_net_1 , \b7_nYhI39s_cry[8] , 
        \b7_nYhI39s_5[8]_net_1 , N_56, G_60_4, N_45, G_60_6, G_60_5, 
        N_76, N_79, \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]_net_1 , N_78, 
        N_81, \b6_Ocm0rW[2] ;
    
    SLE \b3_nUT[0]  (.D(\b6_nUT_IF[0] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  b12_voSc3_gmasbb_RNO (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .Y(
        \b13_nAzGfFM_sLsv3_i_i_0[0] ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[2]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[2]_net_1 ), .Y(\b7_nYhI39s_5[2]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[6]  (.A(
        \b12_uRrc2XfY_rbN[7]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[6]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[6]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[12]  (.D(\b15_uRrc2XfY_rbN_gr[12]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[12]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[11]  (.D(\b12_uRrc2XfY_rbN_5[11]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[11]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[0]  (.D(\status_b2sclk[0] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[0]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  \b13_nAzGfFM_sLsv3_srsts_i_i_a2_0[2]  (
        .A(\b13_nAzGfFM_sLsv3[2]_net_1 ), .B(\b6_nfs_IF[1] ), .C(
        \b3_nfs[4]_net_1 ), .D(b11_PSyil9s_FMZ), .Y(N_56));
    b8_nR_ymqrG_10s_5s_0_0s_0s_1_510_x_0 b11_nUTGT_khWqH (
        .b6_nfs_IF_i_0({\b6_nfs_IF_i_0[1] }), .b6_nUT_IF({
        \b6_nUT_IF[9] , \b6_nUT_IF[8] , \b6_nUT_IF[7] , \b6_nUT_IF[6] , 
        \b6_nUT_IF[5] , \b6_nUT_IF[4] , \b6_nUT_IF[3] , \b6_nUT_IF[2] , 
        \b6_nUT_IF[1] , \b6_nUT_IF[0] }), .b6_nfs_IF({\b6_nfs_IF[4] , 
        \b6_nfs_IF[3] , \b6_nfs_IF[2] , \b6_nfs_IF[1] , \b6_nfs_IF[0] })
        , .IICE_comm2iice_3(IICE_comm2iice[11]), .IICE_comm2iice_0(
        IICE_comm2iice[8]), .IICE_comm2iice_2(IICE_comm2iice[10]), 
        .b4_PLyF(b4_PLyF), .b13_nUTQBgfDb_Z4D(b13_nUTQBgfDb_Z4D), 
        .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), .b16_nYhI39swMeEd_A78(
        b16_nYhI39swMeEd_A78), .b15_nYhI39swMeEd_Mg(
        b15_nYhI39swMeEd_Mg), .b12_vABZ3qsY_Lyh(b12_vABZ3qsY_Lyh), 
        .b11_vABZ3qsY_qH(b11_vABZ3qsY_qH), .b11_vABZ3qsY_XH(
        b11_vABZ3qsY_XH));
    SLE \b3_nUT[6]  (.D(\b6_nUT_IF[6] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[6]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \b6_Ocm0rW_0_0_o2[2]  (.A(
        \b13_nAzGfFM_sLsv3[2]_net_1 ), .B(\b13_nAzGfFM_sLsv3[3]_net_1 )
        , .Y(N_44));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[17]  (.A(
        \b12_uRrc2XfY_rbN[18]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[17]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[17]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[4]  (.D(\b12_uRrc2XfY_rbN_5[4]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[4]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[0]  (.D(\b12_uRrc2XfY_rbN_5[0]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(b12_uRrc2XfY_Lyh));
    SLE \b15_uRrc2XfY_rbN_gs[1]  (.D(\b15_uRrc2XfY_rbN_gr[1]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[10]  (.D(\b15_uRrc2XfY_rbN_gr[10]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[10]_net_1 ));
    SLE \b3_nfs[1]  (.D(\b6_nfs_IF[1] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[5]  (.D(\b15_uRrc2XfY_rbN_gr[5]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \b6_Ocm0rW_0_0[2]  (.A(N_81), .B(
        b13_nAzGfFM_sLsv3_0), .C(N_44), .Y(\b6_Ocm0rW[2] ));
    SLE \b15_uRrc2XfY_rbN_gr[18]  (.D(\b7_nYhI39s[2]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[18]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[14]  (.D(\b12_uRrc2XfY_rbN_5[14]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[14]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIF3AKE[3]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[3]_net_1 ), .D(\b7_nYhI39s_5[3]_net_1 ), .FCI(
        \b7_nYhI39s_cry[2] ), .S(\b7_nYhI39s_s[3] ), .Y(), .FCO(
        \b7_nYhI39s_cry[3] ));
    SLE \b7_nYhI39s[3]  (.D(\b7_nYhI39s_s[3] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[23]  (.D(\b7_nYhI39s[7]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[23]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[24]  (.D(\b15_uRrc2XfY_rbN_gr[24]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[24]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[13]  (.D(\b12_uRrc2XfY_rbN_5[13]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[13]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[1]  (.D(N_94_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b13_nAzGfFM_sLsv3_0));
    SLE \b12_uRrc2XfY_rbN[25]  (.D(\b12_uRrc2XfY_rbN_5[25]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[25]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[13]  (.D(N_104_i_0), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[13]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \b13_nAzGfFM_sLsv3_srsts_i_i_o2[2]  (.A(
        \b13_nAzGfFM_sLsv3[2]_net_1 ), .B(b11_PSyil9s_FMZ), .Y(N_45));
    CFG4 #( .INIT(16'hF0F8) )  \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]  (.A(
        \b13_nAzGfFM_sLsv3[2]_net_1 ), .B(b13_nAzGfFM_sLsv3_0), .C(
        N_56), .D(\b6_nfs_IF[1] ), .Y(
        \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[19]  (.D(\b15_uRrc2XfY_rbN_gr[19]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[19]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[23]  (.A(
        \b12_uRrc2XfY_rbN[24]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[23]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[23]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[19]  (.D(\b12_uRrc2XfY_rbN_5[19]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[19]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[24]  (.A(
        \b12_uRrc2XfY_rbN[25]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[24]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[24]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[25]  (.D(\b15_uRrc2XfY_rbN_gr[25]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[25]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[6]  (.D(\b12_uRrc2XfY_rbN_5[6]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[6]_net_1 ));
    SLE \b3_nUT[1]  (.D(\b6_nUT_IF[1] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[17]  (.D(\b15_uRrc2XfY_rbN_gr[17]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[17]_net_1 ));
    CFG4 #( .INIT(16'h0A0E) )  \b13_nAzGfFM_sLsv3_RNO[4]  (.A(
        \b13_nAzGfFM_sLsv3[4]_net_1 ), .B(b10_nYhI3_umjB_net_1), .C(
        \b6_nfs_IF[1] ), .D(N_79), .Y(N_26_i_0));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNI7BTMQ[7]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[7]_net_1 ), .D(\b7_nYhI39s_5[7]_net_1 ), .FCI(
        \b7_nYhI39s_cry[6] ), .S(\b7_nYhI39s_s[7] ), .Y(), .FCO(
        \b7_nYhI39s_cry[7] ));
    SLE \b7_nYhI39s[6]  (.D(\b7_nYhI39s_s[6] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[6]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[6]  (.D(\b15_uRrc2XfY_rbN_gr[6]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[6]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[14]  (.D(\b15_uRrc2XfY_rbN_gr[14]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[14]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[8]  (.D(\b12_uRrc2XfY_rbN_5[8]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[8]_net_1 ));
    CFG3 #( .INIT(8'hE0) )  un1_b12_uRrc2XfY_rbN10_i (.A(
        IICE_comm2iice[10]), .B(IICE_comm2iice[9]), .C(b11_uRrc2XfY_XH)
        , .Y(un1_b12_uRrc2XfY_rbN10_i_0));
    SLE \b7_nYhI39s[5]  (.D(\b7_nYhI39s_s[5] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[5]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[1]  (.D(\b12_uRrc2XfY_rbN_5[1]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[3]  (.D(\status_b2sclk[3] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[3]_net_1 ));
    SLE \b3_nUT[3]  (.D(\b6_nUT_IF[3] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[15]  (.D(\b15_uRrc2XfY_rbN_gr[15]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[15]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[22]  (.D(\b7_nYhI39s[6]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[22]_net_1 ));
    CFG3 #( .INIT(8'hDF) )  b10_nYhI3_umjB_RNO_0 (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .B(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .C(N_38), .Y(
        un1_b13_nAzGfFM_sLsv3_1_i_0));
    SLE \b3_nfs[0]  (.D(\b6_nfs_IF[0] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[0]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[22]  (.A(
        \b12_uRrc2XfY_rbN[23]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[22]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[22]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[1]  (.A(
        \b12_uRrc2XfY_rbN[2]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[1]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[1]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3_i[0]  (.D(\b6_nfs_IF_i_0[1] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \b15_uRrc2XfY_rbN_gr_RNO[11]  (.A(
        \b13_nAzGfFM_sLsv3[5]_net_1 ), .B(\b13_nAzGfFM_sLsv3[3]_net_1 )
        , .C(b13_nAzGfFM_sLsv3_0), .Y(N_103_i_0));
    CFG4 #( .INIT(16'h0100) )  b10_nYhI3_umjB_RNO_3 (.A(
        \b7_nYhI39s[9]_net_1 ), .B(\b7_nYhI39s[6]_net_1 ), .C(
        \b7_nYhI39s[5]_net_1 ), .D(\b7_nYhI39s[0]_net_1 ), .Y(G_60_5));
    CFG2 #( .INIT(4'h1) )  b10_nYhI3_umjB_RNO_1 (.A(
        \b7_nYhI39s[2]_net_1 ), .B(\b7_nYhI39s[4]_net_1 ), .Y(G_60_4));
    SLE \b15_uRrc2XfY_rbN_gr[12]  (.D(N_44), .CLK(IICE_comm2iice[11]), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b15_uRrc2XfY_rbN_gr[12]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[2]  (.A(
        \b12_uRrc2XfY_rbN[3]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[2]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[9]  (.D(\b15_uRrc2XfY_rbN_gr[9]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[9]_net_1 ));
    SLE \b7_nYhI39s[4]  (.D(\b7_nYhI39s_s[4] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[4]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[8]  (.A(
        \b12_uRrc2XfY_rbN[9]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[8]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[8]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[20]  (.D(\b7_nYhI39s[4]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[20]_net_1 ));
    ARI1 #( .INIT(20'h40E00) )  \b13_nAzGfFM_sLsv3_RNINSNH2[3]  (.A(
        VCC_net_1), .B(N_38), .C(b10_nYhI3_umjB_net_1), .D(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .FCI(VCC_net_1), .S(), .Y(
        \b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .FCO(b7_nYhI39s_cry_cy));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[5]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[5]_net_1 ), .Y(\b7_nYhI39s_5[5]_net_1 ));
    SLE \b7_nYhI39s[9]  (.D(\b7_nYhI39s_s[9] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[9]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \b3_nfs_RNIPR5A1[2]  (.A(\b3_nfs[2]_net_1 )
        , .B(\b3_nfs[4]_net_1 ), .C(\b3_nfs[3]_net_1 ), .Y(N_76));
    SLE \b12_uRrc2XfY_rbN[15]  (.D(\b12_uRrc2XfY_rbN_5[15]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[15]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[11]  (.A(
        \b12_uRrc2XfY_rbN[12]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[11]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[11]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \b13_nAzGfFM_sLsv3_RNO[5]  (.A(
        \b13_nAzGfFM_sLsv3[5]_net_1 ), .B(\b3_nfs[4]_net_1 ), .C(N_45), 
        .D(\b6_nfs_IF[1] ), .Y(N_28_i_0));
    SLE \b15_uRrc2XfY_rbN_gr[10]  (.D(\b6_nfs_IF[4] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[10]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \b13_nAzGfFM_sLsv3_srsts_i_0_a2_1[1]  (.A(
        b8_vABZ3qsY_net_1), .B(\b3_nfs[0]_net_1 ), .C(N_78), .Y(N_81));
    CFG3 #( .INIT(8'h07) )  \b13_nAzGfFM_sLsv3_srsts_i_0_a2[3]  (.A(
        b11_PSyil9s_FMZ), .B(\b13_nAzGfFM_sLsv3[2]_net_1 ), .C(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .Y(N_79));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNI7JJLK[5]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[5]_net_1 ), .D(\b7_nYhI39s_5[5]_net_1 ), .FCI(
        \b7_nYhI39s_cry[4] ), .S(\b7_nYhI39s_s[5] ), .Y(), .FCO(
        \b7_nYhI39s_cry[5] ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[15]  (.A(
        \b12_uRrc2XfY_rbN[16]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[15]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[15]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[10]  (.A(
        \b12_uRrc2XfY_rbN[11]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[10]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[10]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[0]  (.A(
        \b12_uRrc2XfY_rbN[1]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[0]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[0]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[6]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[6]_net_1 ), .Y(\b7_nYhI39s_5[6]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[5]  (.D(N_28_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[5]_net_1 ));
    CFG4 #( .INIT(16'h5FDF) )  b8_vABZ3qsY_RNIG4T32 (.A(
        b13_nAzGfFM_sLsv3_0), .B(N_76), .C(b8_vABZ3qsY_net_1), .D(
        \b3_nfs[0]_net_1 ), .Y(N_38));
    SLE \b15_uRrc2XfY_rbN_gs[21]  (.D(\b15_uRrc2XfY_rbN_gr[21]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[21]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[0]  (.D(\b15_uRrc2XfY_rbN_gr[0]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[0]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[18]  (.A(
        \b12_uRrc2XfY_rbN[19]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[18]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[18]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[7]  (.D(\b6_nfs_IF[1] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[8]  (.D(\b15_uRrc2XfY_rbN_gr[8]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[8]_net_1 ));
    clock2_en_reg_en_5s_x_0 iclksync (.IICE_comm2iice({
        IICE_comm2iice[11]}), .b6_nfs_IF_i_0({\b6_nfs_IF_i_0[1] }), 
        .status_b2sclk({\status_b2sclk[3] , \status_b2sclk[2] , 
        \status_b2sclk[1] , \status_b2sclk[0] }), .b6_nfs_IF({
        \b6_nfs_IF[1] }), .b6_Ocm0rW({\b6_Ocm0rW[2] }), 
        .b13_nAzGfFM_sLsv3_3(\b13_nAzGfFM_sLsv3[5]_net_1 ), 
        .b13_nAzGfFM_sLsv3_0(\b13_nAzGfFM_sLsv3[2]_net_1 ), 
        .b13_nAzGfFM_sLsv3_2(\b13_nAzGfFM_sLsv3[4]_net_1 ), .BW_clk_c(
        BW_clk_c), .N_38(N_38), .N_78(N_78));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIAAINT[8]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[8]_net_1 ), .D(\b7_nYhI39s_5[8]_net_1 ), .FCI(
        \b7_nYhI39s_cry[7] ), .S(\b7_nYhI39s_s[8] ), .Y(), .FCO(
        \b7_nYhI39s_cry[8] ));
    SLE b12_voSc3_gmasbb (.D(\b13_nAzGfFM_sLsv3_i_i_0[0] ), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b8_SoWGfWYY));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[7]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[7]_net_1 ), .Y(\b7_nYhI39s_5[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[6]  (.D(\b6_nfs_IF[0] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[6]_net_1 ));
    SLE \b3_nUT[9]  (.D(\b6_nUT_IF[9] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[9]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[19]  (.D(\b7_nYhI39s[3]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[19]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \b6_Ocm0rW_0_i_a2_1[1]  (.A(
        b10_nYhI3_umjB_net_1), .B(N_76), .C(\b3_nfs[1]_net_1 ), .Y(
        N_78));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[8]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[8]_net_1 ), .Y(\b7_nYhI39s_5[8]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[4]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[4]_net_1 ), .Y(\b7_nYhI39s_5[4]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[24]  (.D(\b7_nYhI39s[8]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[24]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[9]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[9]_net_1 ), .Y(\b7_nYhI39s_5[9]_net_1 ));
    SLE \b7_nYhI39s[0]  (.D(\b7_nYhI39s_s[0] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[0]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[5]  (.D(\b12_uRrc2XfY_rbN_5[5]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[5]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[18]  (.D(\b12_uRrc2XfY_rbN_5[18]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[18]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[16]  (.D(\b15_uRrc2XfY_rbN_gr[16]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[16]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[7]  (.A(
        \b12_uRrc2XfY_rbN[8]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[7]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[7]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[3]  (.D(\b12_uRrc2XfY_rbN_5[3]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[17]  (.D(\b7_nYhI39s[1]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[17]_net_1 ));
    SLE \b7_nYhI39s[2]  (.D(\b7_nYhI39s_s[2] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[2]  (.D(\b15_uRrc2XfY_rbN_gr[2]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[2]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \b15_uRrc2XfY_rbN_gr_RNO[13]  (.A(
        \b13_nAzGfFM_sLsv3[4]_net_1 ), .B(\b13_nAzGfFM_sLsv3[5]_net_1 )
        , .Y(N_104_i_0));
    SLE \b7_nYhI39s[8]  (.D(\b7_nYhI39s_s[8] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[8]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[11]  (.D(\b15_uRrc2XfY_rbN_gr[11]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[11]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[14]  (.D(\b13_nAzGfFM_sLsv3[5]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gr[14]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[3]  (.D(\b15_uRrc2XfY_rbN_gr[3]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[3]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[3]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[3]_net_1 ), .Y(\b7_nYhI39s_5[3]_net_1 ));
    SLE \b3_nUT[5]  (.D(\b6_nUT_IF[5] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[5]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  b10_nYhI3_umjB_RNO (.A(G_60_4), .B(
        G_60_6), .C(G_60_5), .D(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .Y(
        b10_nYhI3_umjB_3));
    SLE \b12_uRrc2XfY_rbN[22]  (.D(\b12_uRrc2XfY_rbN_5[22]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[22]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \b13_nAzGfFM_sLsv3_RNO[3]  (.A(
        b10_nYhI3_umjB_net_1), .B(\b6_nfs_IF[1] ), .C(N_79), .Y(
        N_90_i_0));
    SLE \b3_nfs[4]  (.D(\b6_nfs_IF[4] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[4]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[8]  (.D(\b6_nfs_IF[2] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[8]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[3]  (.A(
        \b12_uRrc2XfY_rbN[4]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[3]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[3]_net_1 ));
    SLE \b3_nfs[2]  (.D(\b6_nfs_IF[2] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[25]  (.D(\b7_nYhI39s[9]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[25]_net_1 ));
    SLE \b3_nUT[8]  (.D(\b6_nUT_IF[8] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[8]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[20]  (.D(\b12_uRrc2XfY_rbN_5[20]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[20]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[9]  (.D(\b12_uRrc2XfY_rbN_5[9]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[9]_net_1 ));
    CFG1 #( .INIT(2'h1) )  b12_voSc3_gmasbb_RNIALH6 (.A(b8_SoWGfWYY), 
        .Y(b8_SoWGfWYY_i));
    SLE \b15_uRrc2XfY_rbN_gs[23]  (.D(\b15_uRrc2XfY_rbN_gr[23]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[23]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[16]  (.A(
        \b12_uRrc2XfY_rbN[17]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[16]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[16]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[15]  (.D(b11_vABZ3qsY_qH), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[15]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[4]  (.D(N_26_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[4]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[2]  (.D(\b12_uRrc2XfY_rbN_5[2]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[2]_net_1 ));
    CFG4 #( .INIT(16'h1311) )  \b13_nAzGfFM_sLsv3_RNO[1]  (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .B(\b6_nfs_IF[1] ), .C(N_81), 
        .D(b13_nAzGfFM_sLsv3_0), .Y(N_94_i_0));
    SLE \b3_nUT[7]  (.D(\b6_nUT_IF[7] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[18]  (.D(\b15_uRrc2XfY_rbN_gr[18]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[18]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[19]  (.A(
        \b12_uRrc2XfY_rbN[20]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[19]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[19]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[21]  (.D(\b12_uRrc2XfY_rbN_5[21]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[21]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[13]  (.A(
        \b12_uRrc2XfY_rbN[14]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[13]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[13]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[14]  (.A(
        \b12_uRrc2XfY_rbN[15]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[14]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[14]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIABCI5[0]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[0]_net_1 ), .D(\b7_nYhI39s_5[0]_net_1 ), .FCI(
        b7_nYhI39s_cry_cy), .S(\b7_nYhI39s_s[0] ), .Y(), .FCO(
        \b7_nYhI39s_cry[0] ));
    SLE \b15_uRrc2XfY_rbN_gs[13]  (.D(\b15_uRrc2XfY_rbN_gr[13]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[13]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  b10_nYhI3_umjB_RNO_2 (.A(
        \b7_nYhI39s[8]_net_1 ), .B(\b7_nYhI39s[7]_net_1 ), .C(
        \b7_nYhI39s[3]_net_1 ), .D(\b7_nYhI39s[1]_net_1 ), .Y(G_60_6));
    CFG4 #( .INIT(16'h1D3F) )  \b13_nAzGfFM_sLsv3_i_RNIST5R2[0]  (.A(
        \b13_nAzGfFM_sLsv3_i[0]_net_1 ), .B(
        \b13_nAzGfFM_sLsv3[3]_net_1 ), .C(b10_nYhI3_umjB_net_1), .D(
        N_38), .Y(N_23_i_0));
    SLE \b12_uRrc2XfY_rbN[16]  (.D(\b12_uRrc2XfY_rbN_5[16]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[16]_net_1 ));
    SLE b10_nYhI3_umjB (.D(b10_nYhI3_umjB_3), .CLK(BW_clk_c), .EN(
        un1_b13_nAzGfFM_sLsv3_1_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b10_nYhI3_umjB_net_1));
    CFG3 #( .INIT(8'h20) )  \b7_nYhI39s_5[0]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[0]_net_1 ), .Y(\b7_nYhI39s_5[0]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[1]  (.D(\status_b2sclk[1] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[1]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[5]  (.A(
        \b12_uRrc2XfY_rbN[6]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[5]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[5]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIAQUKH[4]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[4]_net_1 ), .D(\b7_nYhI39s_5[4]_net_1 ), .FCI(
        \b7_nYhI39s_cry[3] ), .S(\b7_nYhI39s_s[4] ), .Y(), .FCO(
        \b7_nYhI39s_cry[4] ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIMELJB[2]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[2]_net_1 ), .D(\b7_nYhI39s_5[2]_net_1 ), .FCI(
        \b7_nYhI39s_cry[1] ), .S(\b7_nYhI39s_s[2] ), .Y(), .FCO(
        \b7_nYhI39s_cry[2] ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNIVR0J8[1]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[1]_net_1 ), .D(\b7_nYhI39s_5[1]_net_1 ), .FCI(
        \b7_nYhI39s_cry[0] ), .S(\b7_nYhI39s_s[1] ), .Y(), .FCO(
        \b7_nYhI39s_cry[1] ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[21]  (.A(
        \b12_uRrc2XfY_rbN[22]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[21]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[21]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[17]  (.D(\b12_uRrc2XfY_rbN_5[17]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[17]_net_1 ));
    SLE b8_vABZ3qsY (.D(b11_vABZ3qsY_qH), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b8_vABZ3qsY_net_1));
    SLE \b12_uRrc2XfY_rbN[24]  (.D(\b12_uRrc2XfY_rbN_5[24]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[24]_net_1 ));
    ARI1 #( .INIT(20'h61B00) )  \b7_nYhI39s_5_RNI6E8MN[6]  (.A(
        VCC_net_1), .B(\b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(
        \b7_nYhI39s[6]_net_1 ), .D(\b7_nYhI39s_5[6]_net_1 ), .FCI(
        \b7_nYhI39s_cry[5] ), .S(\b7_nYhI39s_s[6] ), .Y(), .FCO(
        \b7_nYhI39s_cry[6] ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[9]  (.A(
        \b12_uRrc2XfY_rbN[10]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[9]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[9]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[23]  (.D(\b12_uRrc2XfY_rbN_5[23]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[23]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[22]  (.D(\b15_uRrc2XfY_rbN_gr[22]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[22]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[12]  (.D(\b12_uRrc2XfY_rbN_5[12]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[12]_net_1 ));
    SLE \b13_nAzGfFM_sLsv3[2]  (.D(N_16), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[2]_net_1 ));
    ARI1 #( .INIT(20'h41B00) )  \b7_nYhI39s_RNO[9]  (.A(VCC_net_1), .B(
        \b13_nAzGfFM_sLsv3_RNINSNH2_Y[3] ), .C(\b7_nYhI39s[9]_net_1 ), 
        .D(\b7_nYhI39s_5[9]_net_1 ), .FCI(\b7_nYhI39s_cry[8] ), .S(
        \b7_nYhI39s_s[9] ), .Y(), .FCO());
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[25]  (.A(b4_PLyF), .B(
        IICE_comm2iice[9]), .C(\b15_uRrc2XfY_rbN_gs[25]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[25]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[20]  (.A(
        \b12_uRrc2XfY_rbN[21]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[20]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[20]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \b12_uRrc2XfY_rbN_5[12]  (.A(
        \b12_uRrc2XfY_rbN[13]_net_1 ), .B(IICE_comm2iice[9]), .C(
        \b15_uRrc2XfY_rbN_gs[12]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[12]_net_1 ));
    SLE \b3_nUT[2]  (.D(\b6_nUT_IF[2] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[2]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[10]  (.D(\b12_uRrc2XfY_rbN_5[10]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[10]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[9]  (.D(\b6_nfs_IF[3] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[9]_net_1 ));
    CFG3 #( .INIT(8'hFD) )  \b7_nYhI39s_5[1]  (.A(b10_nYhI3_umjB_net_1)
        , .B(N_38), .C(\b3_nUT[1]_net_1 ), .Y(\b7_nYhI39s_5[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \b12_uRrc2XfY_rbN_5[4]  (.A(
        IICE_comm2iice[9]), .B(\b12_uRrc2XfY_rbN[5]_net_1 ), .Y(
        \b12_uRrc2XfY_rbN_5[4]_net_1 ));
    SLE \b3_nfs[3]  (.D(\b6_nfs_IF[3] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\b3_nfs[3]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[21]  (.D(\b7_nYhI39s[5]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[21]_net_1 ));
    SLE \b12_uRrc2XfY_rbN[7]  (.D(\b12_uRrc2XfY_rbN_5[7]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(un1_b12_uRrc2XfY_rbN10_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_uRrc2XfY_rbN[7]_net_1 ));
    CFG4 #( .INIT(16'hAAEA) )  \b13_nAzGfFM_sLsv3_srsts_i_i[2]  (.A(
        \b13_nAzGfFM_sLsv3_srsts_i_i_0[2]_net_1 ), .B(N_81), .C(
        b13_nAzGfFM_sLsv3_0), .D(\b6_nfs_IF[1] ), .Y(N_16));
    SLE \b13_nAzGfFM_sLsv3[3]  (.D(N_90_i_0), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_nAzGfFM_sLsv3[3]_net_1 ));
    SLE \b7_nYhI39s[1]  (.D(\b7_nYhI39s_s[1] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[1]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[20]  (.D(\b15_uRrc2XfY_rbN_gr[20]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[20]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[16]  (.D(\b7_nYhI39s[0]_net_1 ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[16]_net_1 ));
    SLE \b7_nYhI39s[7]  (.D(\b7_nYhI39s_s[7] ), .CLK(BW_clk_c), .EN(
        N_23_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b7_nYhI39s[7]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gs[7]  (.D(\b15_uRrc2XfY_rbN_gr[7]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gs[7]_net_1 ));
    SLE \b3_nUT[4]  (.D(\b6_nUT_IF[4] ), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(\b6_nfs_IF_i_0[1] ), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\b3_nUT[4]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[5]  (.D(\b13_nAzGfFM_sLsv3[2]_net_1 ), 
        .CLK(IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b15_uRrc2XfY_rbN_gr[5]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[2]  (.D(\status_b2sclk[2] ), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[2]_net_1 ));
    SLE \b15_uRrc2XfY_rbN_gr[11]  (.D(N_103_i_0), .CLK(
        IICE_comm2iice[11]), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b15_uRrc2XfY_rbN_gr[11]_net_1 ));
    
endmodule


module b3_12m_x(
       b13_nAzGfFM_sLsv3,
       IICE_comm2iice,
       mdiclink_reg,
       b11_OFWNT9L_8tZ,
       b8_SoWGfWYY,
       b8_SoWGfWYY_i,
       BW_clk_c,
       b12_uRrc2XfY_Lyh,
       N_44,
       b11_PSyil9s_FMZ,
       b4_PLyF,
       b11_uRrc2XfY_XH,
       b13_nUTQBgfDb_Z4D,
       b12_nUTQBgfDb_bd,
       b16_nYhI39swMeEd_A78,
       b15_nYhI39swMeEd_Mg,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_XH,
       b7_PSyi3wy,
       b8_PSyiBgYG
    );
output [1:1] b13_nAzGfFM_sLsv3;
input  [11:8] IICE_comm2iice;
input  [154:0] mdiclink_reg;
input  [154:0] b11_OFWNT9L_8tZ;
output b8_SoWGfWYY;
output b8_SoWGfWYY_i;
input  BW_clk_c;
output b12_uRrc2XfY_Lyh;
output N_44;
output b11_PSyil9s_FMZ;
input  b4_PLyF;
input  b11_uRrc2XfY_XH;
output b13_nUTQBgfDb_Z4D;
input  b12_nUTQBgfDb_bd;
output b16_nYhI39swMeEd_A78;
input  b15_nYhI39swMeEd_Mg;
output b12_vABZ3qsY_Lyh;
input  b11_vABZ3qsY_XH;
output b7_PSyi3wy;
input  b8_PSyiBgYG;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    b7_PfFzrNY_x_0 b4_PfFz (.mdiclink_reg({mdiclink_reg[154], 
        mdiclink_reg[153], mdiclink_reg[152], mdiclink_reg[151], 
        mdiclink_reg[150], mdiclink_reg[149], mdiclink_reg[148], 
        mdiclink_reg[147], mdiclink_reg[146], mdiclink_reg[145], 
        mdiclink_reg[144], mdiclink_reg[143], mdiclink_reg[142], 
        mdiclink_reg[141], mdiclink_reg[140], mdiclink_reg[139], 
        mdiclink_reg[138], mdiclink_reg[137], mdiclink_reg[136], 
        mdiclink_reg[135], mdiclink_reg[134], mdiclink_reg[133], 
        mdiclink_reg[132], mdiclink_reg[131], mdiclink_reg[130], 
        mdiclink_reg[129], mdiclink_reg[128], mdiclink_reg[127], 
        mdiclink_reg[126], mdiclink_reg[125], mdiclink_reg[124], 
        mdiclink_reg[123], mdiclink_reg[122], mdiclink_reg[121], 
        mdiclink_reg[120], mdiclink_reg[119], mdiclink_reg[118], 
        mdiclink_reg[117], mdiclink_reg[116], mdiclink_reg[115], 
        mdiclink_reg[114], mdiclink_reg[113], mdiclink_reg[112], 
        mdiclink_reg[111], mdiclink_reg[110], mdiclink_reg[109], 
        mdiclink_reg[108], mdiclink_reg[107], mdiclink_reg[106], 
        mdiclink_reg[105], mdiclink_reg[104], mdiclink_reg[103], 
        mdiclink_reg[102], mdiclink_reg[101], mdiclink_reg[100], 
        mdiclink_reg[99], mdiclink_reg[98], mdiclink_reg[97], 
        mdiclink_reg[96], mdiclink_reg[95], mdiclink_reg[94], 
        mdiclink_reg[93], mdiclink_reg[92], mdiclink_reg[91], 
        mdiclink_reg[90], mdiclink_reg[89], mdiclink_reg[88], 
        mdiclink_reg[87], mdiclink_reg[86], mdiclink_reg[85], 
        mdiclink_reg[84], mdiclink_reg[83], mdiclink_reg[82], 
        mdiclink_reg[81], mdiclink_reg[80], mdiclink_reg[79], 
        mdiclink_reg[78], mdiclink_reg[77], mdiclink_reg[76], 
        mdiclink_reg[75], mdiclink_reg[74], mdiclink_reg[73], 
        mdiclink_reg[72], mdiclink_reg[71], mdiclink_reg[70], 
        mdiclink_reg[69], mdiclink_reg[68], mdiclink_reg[67], 
        mdiclink_reg[66], mdiclink_reg[65], mdiclink_reg[64], 
        mdiclink_reg[63], mdiclink_reg[62], mdiclink_reg[61], 
        mdiclink_reg[60], mdiclink_reg[59], mdiclink_reg[58], 
        mdiclink_reg[57], mdiclink_reg[56], mdiclink_reg[55], 
        mdiclink_reg[54], mdiclink_reg[53], mdiclink_reg[52], 
        mdiclink_reg[51], mdiclink_reg[50], mdiclink_reg[49], 
        mdiclink_reg[48], mdiclink_reg[47], mdiclink_reg[46], 
        mdiclink_reg[45], mdiclink_reg[44], mdiclink_reg[43], 
        mdiclink_reg[42], mdiclink_reg[41], mdiclink_reg[40], 
        mdiclink_reg[39], mdiclink_reg[38], mdiclink_reg[37], 
        mdiclink_reg[36], mdiclink_reg[35], mdiclink_reg[34], 
        mdiclink_reg[33], mdiclink_reg[32], mdiclink_reg[31], 
        mdiclink_reg[30], mdiclink_reg[29], mdiclink_reg[28], 
        mdiclink_reg[27], mdiclink_reg[26], mdiclink_reg[25], 
        mdiclink_reg[24], mdiclink_reg[23], mdiclink_reg[22], 
        mdiclink_reg[21], mdiclink_reg[20], mdiclink_reg[19], 
        mdiclink_reg[18], mdiclink_reg[17], mdiclink_reg[16], 
        mdiclink_reg[15], mdiclink_reg[14], mdiclink_reg[13], 
        mdiclink_reg[12], mdiclink_reg[11], mdiclink_reg[10], 
        mdiclink_reg[9], mdiclink_reg[8], mdiclink_reg[7], 
        mdiclink_reg[6], mdiclink_reg[5], mdiclink_reg[4], 
        mdiclink_reg[3], mdiclink_reg[2], mdiclink_reg[1], 
        mdiclink_reg[0]}), .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[154], 
        b11_OFWNT9L_8tZ[153], b11_OFWNT9L_8tZ[152], 
        b11_OFWNT9L_8tZ[151], b11_OFWNT9L_8tZ[150], 
        b11_OFWNT9L_8tZ[149], b11_OFWNT9L_8tZ[148], 
        b11_OFWNT9L_8tZ[147], b11_OFWNT9L_8tZ[146], 
        b11_OFWNT9L_8tZ[145], b11_OFWNT9L_8tZ[144], 
        b11_OFWNT9L_8tZ[143], b11_OFWNT9L_8tZ[142], 
        b11_OFWNT9L_8tZ[141], b11_OFWNT9L_8tZ[140], 
        b11_OFWNT9L_8tZ[139], b11_OFWNT9L_8tZ[138], 
        b11_OFWNT9L_8tZ[137], b11_OFWNT9L_8tZ[136], 
        b11_OFWNT9L_8tZ[135], b11_OFWNT9L_8tZ[134], 
        b11_OFWNT9L_8tZ[133], b11_OFWNT9L_8tZ[132], 
        b11_OFWNT9L_8tZ[131], b11_OFWNT9L_8tZ[130], 
        b11_OFWNT9L_8tZ[129], b11_OFWNT9L_8tZ[128], 
        b11_OFWNT9L_8tZ[127], b11_OFWNT9L_8tZ[126], 
        b11_OFWNT9L_8tZ[125], b11_OFWNT9L_8tZ[124], 
        b11_OFWNT9L_8tZ[123], b11_OFWNT9L_8tZ[122], 
        b11_OFWNT9L_8tZ[121], b11_OFWNT9L_8tZ[120], 
        b11_OFWNT9L_8tZ[119], b11_OFWNT9L_8tZ[118], 
        b11_OFWNT9L_8tZ[117], b11_OFWNT9L_8tZ[116], 
        b11_OFWNT9L_8tZ[115], b11_OFWNT9L_8tZ[114], 
        b11_OFWNT9L_8tZ[113], b11_OFWNT9L_8tZ[112], 
        b11_OFWNT9L_8tZ[111], b11_OFWNT9L_8tZ[110], 
        b11_OFWNT9L_8tZ[109], b11_OFWNT9L_8tZ[108], 
        b11_OFWNT9L_8tZ[107], b11_OFWNT9L_8tZ[106], 
        b11_OFWNT9L_8tZ[105], b11_OFWNT9L_8tZ[104], 
        b11_OFWNT9L_8tZ[103], b11_OFWNT9L_8tZ[102], 
        b11_OFWNT9L_8tZ[101], b11_OFWNT9L_8tZ[100], 
        b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], b11_OFWNT9L_8tZ[97], 
        b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], b11_OFWNT9L_8tZ[94], 
        b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], b11_OFWNT9L_8tZ[91], 
        b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], b11_OFWNT9L_8tZ[88], 
        b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], b11_OFWNT9L_8tZ[85], 
        b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], b11_OFWNT9L_8tZ[82], 
        b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], b11_OFWNT9L_8tZ[79], 
        b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], b11_OFWNT9L_8tZ[76], 
        b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], b11_OFWNT9L_8tZ[73], 
        b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], b11_OFWNT9L_8tZ[70], 
        b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], b11_OFWNT9L_8tZ[67], 
        b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], b11_OFWNT9L_8tZ[64], 
        b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], b11_OFWNT9L_8tZ[61], 
        b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], b11_OFWNT9L_8tZ[58], 
        b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], b11_OFWNT9L_8tZ[55], 
        b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], b11_OFWNT9L_8tZ[52], 
        b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], b11_OFWNT9L_8tZ[49], 
        b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], b11_OFWNT9L_8tZ[46], 
        b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], b11_OFWNT9L_8tZ[43], 
        b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], b11_OFWNT9L_8tZ[40], 
        b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], b11_OFWNT9L_8tZ[37], 
        b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], b11_OFWNT9L_8tZ[34], 
        b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], b11_OFWNT9L_8tZ[31], 
        b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], b11_OFWNT9L_8tZ[28], 
        b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], b11_OFWNT9L_8tZ[25], 
        b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], b11_OFWNT9L_8tZ[22], 
        b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], b11_OFWNT9L_8tZ[19], 
        b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], b11_OFWNT9L_8tZ[16], 
        b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], b11_OFWNT9L_8tZ[13], 
        b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], b11_OFWNT9L_8tZ[10], 
        b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], b11_OFWNT9L_8tZ[7], 
        b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], b11_OFWNT9L_8tZ[4], 
        b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], b11_OFWNT9L_8tZ[1], 
        b11_OFWNT9L_8tZ[0]}), .IICE_comm2iice({IICE_comm2iice[11], 
        IICE_comm2iice[10]}), .b11_PSyil9s_FMZ(b11_PSyil9s_FMZ), 
        .BW_clk_c(BW_clk_c), .b7_PSyi3wy(b7_PSyi3wy), .b4_PLyF(b4_PLyF)
        , .b8_PSyiBgYG(b8_PSyiBgYG));
    GND GND (.Y(GND_net_1));
    b7_OCByLXC_Z1_x_0 b5_nUTGT (.IICE_comm2iice({IICE_comm2iice[11], 
        IICE_comm2iice[10], IICE_comm2iice[9], IICE_comm2iice[8]}), 
        .b13_nAzGfFM_sLsv3_0(b13_nAzGfFM_sLsv3[1]), .b8_SoWGfWYY(
        b8_SoWGfWYY), .b8_SoWGfWYY_i(b8_SoWGfWYY_i), .BW_clk_c(
        BW_clk_c), .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh), .N_44(N_44), 
        .b11_PSyil9s_FMZ(b11_PSyil9s_FMZ), .b4_PLyF(b4_PLyF), 
        .b11_uRrc2XfY_XH(b11_uRrc2XfY_XH), .b13_nUTQBgfDb_Z4D(
        b13_nUTQBgfDb_Z4D), .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), 
        .b16_nYhI39swMeEd_A78(b16_nYhI39swMeEd_A78), 
        .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), .b12_vABZ3qsY_Lyh(
        b12_vABZ3qsY_Lyh), .b11_vABZ3qsY_XH(b11_vABZ3qsY_XH));
    
endmodule


module b13_vFW_xNywD_EdR_161s_10s_1024s_0s_x_0(
       IICE_comm2iice,
       b12_2_St6KCa_jHv,
       b7_vFW_PlM,
       b11_OFWNT9L_8tZ,
       b9_v_mzCDYXs_2,
       b9_v_mzCDYXs_1,
       b9_v_mzCDYXs_0,
       b9_v_mzCDYXs,
       b9_v_mzCDYXs_8,
       b9_v_mzCDYXs_7,
       b9_v_mzCDYXs_6,
       b9_v_mzCDYXs_5,
       b9_v_mzCDYXs_4,
       b9_v_mzCDYXs_3,
       BW_clk_c,
       b4_2o_z
    );
input  [11:11] IICE_comm2iice;
input  [9:0] b12_2_St6KCa_jHv;
output [154:0] b7_vFW_PlM;
input  [154:0] b11_OFWNT9L_8tZ;
input  b9_v_mzCDYXs_2;
input  b9_v_mzCDYXs_1;
input  b9_v_mzCDYXs_0;
input  b9_v_mzCDYXs;
input  b9_v_mzCDYXs_8;
input  b9_v_mzCDYXs_7;
input  b9_v_mzCDYXs_6;
input  b9_v_mzCDYXs_5;
input  b9_v_mzCDYXs_4;
input  b9_v_mzCDYXs_3;
input  BW_clk_c;
input  b4_2o_z;

    wire VCC_net_1, GND_net_1;
    
    RAM1K18 b3_SoW_b3_SoW_0_1 (.A_DOUT({b7_vFW_PlM[35], b7_vFW_PlM[34], 
        b7_vFW_PlM[33], b7_vFW_PlM[32], b7_vFW_PlM[31], b7_vFW_PlM[30], 
        b7_vFW_PlM[29], b7_vFW_PlM[28], b7_vFW_PlM[27], b7_vFW_PlM[26], 
        b7_vFW_PlM[25], b7_vFW_PlM[24], b7_vFW_PlM[23], b7_vFW_PlM[22], 
        b7_vFW_PlM[21], b7_vFW_PlM[20], b7_vFW_PlM[19], b7_vFW_PlM[18]})
        , .B_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, 
        nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17}), .BUSY(), 
        .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[35], b11_OFWNT9L_8tZ[34], b11_OFWNT9L_8tZ[33], 
        b11_OFWNT9L_8tZ[32], b11_OFWNT9L_8tZ[31], b11_OFWNT9L_8tZ[30], 
        b11_OFWNT9L_8tZ[29], b11_OFWNT9L_8tZ[28], b11_OFWNT9L_8tZ[27], 
        b11_OFWNT9L_8tZ[26], b11_OFWNT9L_8tZ[25], b11_OFWNT9L_8tZ[24], 
        b11_OFWNT9L_8tZ[23], b11_OFWNT9L_8tZ[22], b11_OFWNT9L_8tZ[21], 
        b11_OFWNT9L_8tZ[20], b11_OFWNT9L_8tZ[19], b11_OFWNT9L_8tZ[18]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_0 (.A_DOUT({b7_vFW_PlM[17], b7_vFW_PlM[16], 
        b7_vFW_PlM[15], b7_vFW_PlM[14], b7_vFW_PlM[13], b7_vFW_PlM[12], 
        b7_vFW_PlM[11], b7_vFW_PlM[10], b7_vFW_PlM[9], b7_vFW_PlM[8], 
        b7_vFW_PlM[7], b7_vFW_PlM[6], b7_vFW_PlM[5], b7_vFW_PlM[4], 
        b7_vFW_PlM[3], b7_vFW_PlM[2], b7_vFW_PlM[1], b7_vFW_PlM[0]}), 
        .B_DOUT({nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, nc26, 
        nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35}), .BUSY()
        , .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[17], b11_OFWNT9L_8tZ[16], b11_OFWNT9L_8tZ[15], 
        b11_OFWNT9L_8tZ[14], b11_OFWNT9L_8tZ[13], b11_OFWNT9L_8tZ[12], 
        b11_OFWNT9L_8tZ[11], b11_OFWNT9L_8tZ[10], b11_OFWNT9L_8tZ[9], 
        b11_OFWNT9L_8tZ[8], b11_OFWNT9L_8tZ[7], b11_OFWNT9L_8tZ[6], 
        b11_OFWNT9L_8tZ[5], b11_OFWNT9L_8tZ[4], b11_OFWNT9L_8tZ[3], 
        b11_OFWNT9L_8tZ[2], b11_OFWNT9L_8tZ[1], b11_OFWNT9L_8tZ[0]}), 
        .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    GND GND (.Y(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_4 (.A_DOUT({b7_vFW_PlM[89], b7_vFW_PlM[88], 
        b7_vFW_PlM[87], b7_vFW_PlM[86], b7_vFW_PlM[85], b7_vFW_PlM[84], 
        b7_vFW_PlM[83], b7_vFW_PlM[82], b7_vFW_PlM[81], b7_vFW_PlM[80], 
        b7_vFW_PlM[79], b7_vFW_PlM[78], b7_vFW_PlM[77], b7_vFW_PlM[76], 
        b7_vFW_PlM[75], b7_vFW_PlM[74], b7_vFW_PlM[73], b7_vFW_PlM[72]})
        , .B_DOUT({nc36, nc37, nc38, nc39, nc40, nc41, nc42, nc43, 
        nc44, nc45, nc46, nc47, nc48, nc49, nc50, nc51, nc52, nc53}), 
        .BUSY(), .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(
        IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), 
        .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[89], b11_OFWNT9L_8tZ[88], b11_OFWNT9L_8tZ[87], 
        b11_OFWNT9L_8tZ[86], b11_OFWNT9L_8tZ[85], b11_OFWNT9L_8tZ[84], 
        b11_OFWNT9L_8tZ[83], b11_OFWNT9L_8tZ[82], b11_OFWNT9L_8tZ[81], 
        b11_OFWNT9L_8tZ[80], b11_OFWNT9L_8tZ[79], b11_OFWNT9L_8tZ[78], 
        b11_OFWNT9L_8tZ[77], b11_OFWNT9L_8tZ[76], b11_OFWNT9L_8tZ[75], 
        b11_OFWNT9L_8tZ[74], b11_OFWNT9L_8tZ[73], b11_OFWNT9L_8tZ[72]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_7 (.A_DOUT({b7_vFW_PlM[143], 
        b7_vFW_PlM[142], b7_vFW_PlM[141], b7_vFW_PlM[140], 
        b7_vFW_PlM[139], b7_vFW_PlM[138], b7_vFW_PlM[137], 
        b7_vFW_PlM[136], b7_vFW_PlM[135], b7_vFW_PlM[134], 
        b7_vFW_PlM[133], b7_vFW_PlM[132], b7_vFW_PlM[131], 
        b7_vFW_PlM[130], b7_vFW_PlM[129], b7_vFW_PlM[128], 
        b7_vFW_PlM[127], b7_vFW_PlM[126]}), .B_DOUT({nc54, nc55, nc56, 
        nc57, nc58, nc59, nc60, nc61, nc62, nc63, nc64, nc65, nc66, 
        nc67, nc68, nc69, nc70, nc71}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[143], b11_OFWNT9L_8tZ[142], 
        b11_OFWNT9L_8tZ[141], b11_OFWNT9L_8tZ[140], 
        b11_OFWNT9L_8tZ[139], b11_OFWNT9L_8tZ[138], 
        b11_OFWNT9L_8tZ[137], b11_OFWNT9L_8tZ[136], 
        b11_OFWNT9L_8tZ[135], b11_OFWNT9L_8tZ[134], 
        b11_OFWNT9L_8tZ[133], b11_OFWNT9L_8tZ[132], 
        b11_OFWNT9L_8tZ[131], b11_OFWNT9L_8tZ[130], 
        b11_OFWNT9L_8tZ[129], b11_OFWNT9L_8tZ[128], 
        b11_OFWNT9L_8tZ[127], b11_OFWNT9L_8tZ[126]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_6 (.A_DOUT({b7_vFW_PlM[125], 
        b7_vFW_PlM[124], b7_vFW_PlM[123], b7_vFW_PlM[122], 
        b7_vFW_PlM[121], b7_vFW_PlM[120], b7_vFW_PlM[119], 
        b7_vFW_PlM[118], b7_vFW_PlM[117], b7_vFW_PlM[116], 
        b7_vFW_PlM[115], b7_vFW_PlM[114], b7_vFW_PlM[113], 
        b7_vFW_PlM[112], b7_vFW_PlM[111], b7_vFW_PlM[110], 
        b7_vFW_PlM[109], b7_vFW_PlM[108]}), .B_DOUT({nc72, nc73, nc74, 
        nc75, nc76, nc77, nc78, nc79, nc80, nc81, nc82, nc83, nc84, 
        nc85, nc86, nc87, nc88, nc89}), .BUSY(), .A_CLK(
        IICE_comm2iice[11]), .A_DOUT_CLK(IICE_comm2iice[11]), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, b9_v_mzCDYXs_4, 
        b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, b9_v_mzCDYXs_8, 
        b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, b9_v_mzCDYXs_2, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[125], b11_OFWNT9L_8tZ[124], 
        b11_OFWNT9L_8tZ[123], b11_OFWNT9L_8tZ[122], 
        b11_OFWNT9L_8tZ[121], b11_OFWNT9L_8tZ[120], 
        b11_OFWNT9L_8tZ[119], b11_OFWNT9L_8tZ[118], 
        b11_OFWNT9L_8tZ[117], b11_OFWNT9L_8tZ[116], 
        b11_OFWNT9L_8tZ[115], b11_OFWNT9L_8tZ[114], 
        b11_OFWNT9L_8tZ[113], b11_OFWNT9L_8tZ[112], 
        b11_OFWNT9L_8tZ[111], b11_OFWNT9L_8tZ[110], 
        b11_OFWNT9L_8tZ[109], b11_OFWNT9L_8tZ[108]}), .B_ADDR({
        b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], 
        b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], 
        b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], 
        b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_5 (.A_DOUT({b7_vFW_PlM[107], 
        b7_vFW_PlM[106], b7_vFW_PlM[105], b7_vFW_PlM[104], 
        b7_vFW_PlM[103], b7_vFW_PlM[102], b7_vFW_PlM[101], 
        b7_vFW_PlM[100], b7_vFW_PlM[99], b7_vFW_PlM[98], 
        b7_vFW_PlM[97], b7_vFW_PlM[96], b7_vFW_PlM[95], b7_vFW_PlM[94], 
        b7_vFW_PlM[93], b7_vFW_PlM[92], b7_vFW_PlM[91], b7_vFW_PlM[90]})
        , .B_DOUT({nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97, 
        nc98, nc99, nc100, nc101, nc102, nc103, nc104, nc105, nc106, 
        nc107}), .BUSY(), .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(
        IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), 
        .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[107], b11_OFWNT9L_8tZ[106], 
        b11_OFWNT9L_8tZ[105], b11_OFWNT9L_8tZ[104], 
        b11_OFWNT9L_8tZ[103], b11_OFWNT9L_8tZ[102], 
        b11_OFWNT9L_8tZ[101], b11_OFWNT9L_8tZ[100], 
        b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], b11_OFWNT9L_8tZ[97], 
        b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], b11_OFWNT9L_8tZ[94], 
        b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], b11_OFWNT9L_8tZ[91], 
        b11_OFWNT9L_8tZ[90]}), .B_ADDR({b12_2_St6KCa_jHv[9], 
        b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], 
        b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], 
        b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, 
        b4_2o_z}), .A_EN(VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({
        VCC_net_1, GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(
        VCC_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(
        GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_3 (.A_DOUT({b7_vFW_PlM[71], b7_vFW_PlM[70], 
        b7_vFW_PlM[69], b7_vFW_PlM[68], b7_vFW_PlM[67], b7_vFW_PlM[66], 
        b7_vFW_PlM[65], b7_vFW_PlM[64], b7_vFW_PlM[63], b7_vFW_PlM[62], 
        b7_vFW_PlM[61], b7_vFW_PlM[60], b7_vFW_PlM[59], b7_vFW_PlM[58], 
        b7_vFW_PlM[57], b7_vFW_PlM[56], b7_vFW_PlM[55], b7_vFW_PlM[54]})
        , .B_DOUT({nc108, nc109, nc110, nc111, nc112, nc113, nc114, 
        nc115, nc116, nc117, nc118, nc119, nc120, nc121, nc122, nc123, 
        nc124, nc125}), .BUSY(), .A_CLK(IICE_comm2iice[11]), 
        .A_DOUT_CLK(IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), 
        .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1})
        , .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[71], b11_OFWNT9L_8tZ[70], b11_OFWNT9L_8tZ[69], 
        b11_OFWNT9L_8tZ[68], b11_OFWNT9L_8tZ[67], b11_OFWNT9L_8tZ[66], 
        b11_OFWNT9L_8tZ[65], b11_OFWNT9L_8tZ[64], b11_OFWNT9L_8tZ[63], 
        b11_OFWNT9L_8tZ[62], b11_OFWNT9L_8tZ[61], b11_OFWNT9L_8tZ[60], 
        b11_OFWNT9L_8tZ[59], b11_OFWNT9L_8tZ[58], b11_OFWNT9L_8tZ[57], 
        b11_OFWNT9L_8tZ[56], b11_OFWNT9L_8tZ[55], b11_OFWNT9L_8tZ[54]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_2 (.A_DOUT({b7_vFW_PlM[53], b7_vFW_PlM[52], 
        b7_vFW_PlM[51], b7_vFW_PlM[50], b7_vFW_PlM[49], b7_vFW_PlM[48], 
        b7_vFW_PlM[47], b7_vFW_PlM[46], b7_vFW_PlM[45], b7_vFW_PlM[44], 
        b7_vFW_PlM[43], b7_vFW_PlM[42], b7_vFW_PlM[41], b7_vFW_PlM[40], 
        b7_vFW_PlM[39], b7_vFW_PlM[38], b7_vFW_PlM[37], b7_vFW_PlM[36]})
        , .B_DOUT({nc126, nc127, nc128, nc129, nc130, nc131, nc132, 
        nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, nc141, 
        nc142, nc143}), .BUSY(), .A_CLK(IICE_comm2iice[11]), 
        .A_DOUT_CLK(IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), 
        .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1})
        , .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        b11_OFWNT9L_8tZ[53], b11_OFWNT9L_8tZ[52], b11_OFWNT9L_8tZ[51], 
        b11_OFWNT9L_8tZ[50], b11_OFWNT9L_8tZ[49], b11_OFWNT9L_8tZ[48], 
        b11_OFWNT9L_8tZ[47], b11_OFWNT9L_8tZ[46], b11_OFWNT9L_8tZ[45], 
        b11_OFWNT9L_8tZ[44], b11_OFWNT9L_8tZ[43], b11_OFWNT9L_8tZ[42], 
        b11_OFWNT9L_8tZ[41], b11_OFWNT9L_8tZ[40], b11_OFWNT9L_8tZ[39], 
        b11_OFWNT9L_8tZ[38], b11_OFWNT9L_8tZ[37], b11_OFWNT9L_8tZ[36]})
        , .B_ADDR({b12_2_St6KCa_jHv[9], b12_2_St6KCa_jHv[8], 
        b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], b12_2_St6KCa_jHv[5], 
        b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], b12_2_St6KCa_jHv[2], 
        b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, b4_2o_z}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(GND_net_1));
    RAM1K18 b3_SoW_b3_SoW_0_8 (.A_DOUT({nc144, nc145, nc146, nc147, 
        nc148, nc149, nc150, b7_vFW_PlM[154], b7_vFW_PlM[153], 
        b7_vFW_PlM[152], b7_vFW_PlM[151], b7_vFW_PlM[150], 
        b7_vFW_PlM[149], b7_vFW_PlM[148], b7_vFW_PlM[147], 
        b7_vFW_PlM[146], b7_vFW_PlM[145], b7_vFW_PlM[144]}), .B_DOUT({
        nc151, nc152, nc153, nc154, nc155, nc156, nc157, nc158, nc159, 
        nc160, nc161, nc162, nc163, nc164, nc165, nc166, nc167, nc168})
        , .BUSY(), .A_CLK(IICE_comm2iice[11]), .A_DOUT_CLK(
        IICE_comm2iice[11]), .A_ARST_N(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), 
        .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({b9_v_mzCDYXs_3, 
        b9_v_mzCDYXs_4, b9_v_mzCDYXs_5, b9_v_mzCDYXs_6, b9_v_mzCDYXs_7, 
        b9_v_mzCDYXs_8, b9_v_mzCDYXs, b9_v_mzCDYXs_0, b9_v_mzCDYXs_1, 
        b9_v_mzCDYXs_2, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({GND_net_1, GND_net_1}), .B_CLK(BW_clk_c), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({VCC_net_1, VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(
        VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, b11_OFWNT9L_8tZ[154], b11_OFWNT9L_8tZ[153], 
        b11_OFWNT9L_8tZ[152], b11_OFWNT9L_8tZ[151], 
        b11_OFWNT9L_8tZ[150], b11_OFWNT9L_8tZ[149], 
        b11_OFWNT9L_8tZ[148], b11_OFWNT9L_8tZ[147], 
        b11_OFWNT9L_8tZ[146], b11_OFWNT9L_8tZ[145], 
        b11_OFWNT9L_8tZ[144]}), .B_ADDR({b12_2_St6KCa_jHv[9], 
        b12_2_St6KCa_jHv[8], b12_2_St6KCa_jHv[7], b12_2_St6KCa_jHv[6], 
        b12_2_St6KCa_jHv[5], b12_2_St6KCa_jHv[4], b12_2_St6KCa_jHv[3], 
        b12_2_St6KCa_jHv[2], b12_2_St6KCa_jHv[1], b12_2_St6KCa_jHv[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .B_WEN({b4_2o_z, 
        b4_2o_z}), .A_EN(VCC_net_1), .A_DOUT_LAT(GND_net_1), .A_WIDTH({
        VCC_net_1, GND_net_1, GND_net_1}), .A_WMODE(VCC_net_1), .B_EN(
        VCC_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, 
        GND_net_1, GND_net_1}), .B_WMODE(VCC_net_1), .SII_LOCK(
        GND_net_1));
    
endmodule


module b19_nczQ_DYg_YFaRM_oUoP_24s_1s_x_0(
       b12_PSyi_KyDbLbb,
       b8_FZFFLXYE,
       IICE_comm2iice_6,
       IICE_comm2iice_4,
       IICE_comm2iice_0,
       ttdo,
       b8_jAA_KlCO,
       un1_b13_PLF_2grFt_FH911_i_a2_0_1,
       un1_b13_PLF_2grFt_FH911_i_a2_0_2,
       N_14_1
    );
input  [9:0] b12_PSyi_KyDbLbb;
input  [9:0] b8_FZFFLXYE;
input  IICE_comm2iice_6;
input  IICE_comm2iice_4;
input  IICE_comm2iice_0;
output ttdo;
input  b8_jAA_KlCO;
input  un1_b13_PLF_2grFt_FH911_i_a2_0_1;
input  un1_b13_PLF_2grFt_FH911_i_a2_0_2;
input  N_14_1;

    wire \b13_PLF_2grFt_FH9[22] , VCC_net_1, 
        \b13_PLF_2grFt_FH9_10[22] , N_14, GND_net_1, 
        \b13_PLF_2grFt_FH9[23] , \b13_PLF_2grFt_FH9_10[23] , 
        \b13_PLF_2grFt_FH9[7] , \b13_PLF_2grFt_FH9_10[7] , 
        \b13_PLF_2grFt_FH9[8] , \b13_PLF_2grFt_FH9_10[8] , 
        \b13_PLF_2grFt_FH9[9] , \b13_PLF_2grFt_FH9_10[9] , 
        \b13_PLF_2grFt_FH9[10] , \b13_PLF_2grFt_FH9_10[10] , 
        \b13_PLF_2grFt_FH9[11] , \b13_PLF_2grFt_FH9_10[11] , 
        \b13_PLF_2grFt_FH9[12] , \b13_PLF_2grFt_FH9_10[12] , 
        \b13_PLF_2grFt_FH9[13] , \b13_PLF_2grFt_FH9_10[13] , 
        \b13_PLF_2grFt_FH9[14] , \b13_PLF_2grFt_FH9_10[14] , 
        \b13_PLF_2grFt_FH9[15] , \b13_PLF_2grFt_FH9_10[15] , 
        \b13_PLF_2grFt_FH9[16] , \b13_PLF_2grFt_FH9_10[16] , 
        \b13_PLF_2grFt_FH9[17] , \b13_PLF_2grFt_FH9_10[17] , 
        \b13_PLF_2grFt_FH9[18] , \b13_PLF_2grFt_FH9_10[18] , 
        \b13_PLF_2grFt_FH9[19] , \b13_PLF_2grFt_FH9_10[19] , 
        \b13_PLF_2grFt_FH9[20] , \b13_PLF_2grFt_FH9_10[20] , 
        \b13_PLF_2grFt_FH9[21] , \b13_PLF_2grFt_FH9_10[21] , 
        \b13_PLF_2grFt_FH9_10[0] , \b13_PLF_2grFt_FH9[1] , 
        \b13_PLF_2grFt_FH9_10[1] , \b13_PLF_2grFt_FH9[2] , 
        \b13_PLF_2grFt_FH9_10[2] , \b13_PLF_2grFt_FH9[3] , 
        \b13_PLF_2grFt_FH9_10[3] , \b13_PLF_2grFt_FH9[4] , 
        \b13_PLF_2grFt_FH9_10[4] , \b13_PLF_2grFt_FH9[5] , 
        \b13_PLF_2grFt_FH9_10[5] , \b13_PLF_2grFt_FH9[6] , 
        \b13_PLF_2grFt_FH9_10[6] ;
    
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_10[0]  (.A(
        IICE_comm2iice_4), .B(\b13_PLF_2grFt_FH9[1] ), .Y(
        \b13_PLF_2grFt_FH9_10[0] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[19]  (.A(
        b12_PSyi_KyDbLbb[5]), .B(\b13_PLF_2grFt_FH9[20] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[19] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[2]  (.D(\b13_PLF_2grFt_FH9_10[2] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[2] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[22]  (.A(
        b12_PSyi_KyDbLbb[8]), .B(\b13_PLF_2grFt_FH9[23] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[22] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[15]  (.A(
        b12_PSyi_KyDbLbb[1]), .B(\b13_PLF_2grFt_FH9[16] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[15] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[2]  (.A(
        b8_jAA_KlCO), .B(\b13_PLF_2grFt_FH9[3] ), .C(IICE_comm2iice_4), 
        .Y(\b13_PLF_2grFt_FH9_10[2] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[5]  (.D(\b13_PLF_2grFt_FH9_10[5] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[5] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[5]  (.A(
        b8_FZFFLXYE[1]), .B(\b13_PLF_2grFt_FH9[6] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[5] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[16]  (.D(\b13_PLF_2grFt_FH9_10[16] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[16] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_10[1]  (.A(
        IICE_comm2iice_4), .B(\b13_PLF_2grFt_FH9[2] ), .Y(
        \b13_PLF_2grFt_FH9_10[1] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_10[3]  (.A(
        IICE_comm2iice_4), .B(\b13_PLF_2grFt_FH9[4] ), .Y(
        \b13_PLF_2grFt_FH9_10[3] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[10]  (.D(\b13_PLF_2grFt_FH9_10[10] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[10] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[12]  (.A(
        b8_FZFFLXYE[8]), .B(\b13_PLF_2grFt_FH9[13] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[12] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[23]  (.D(\b13_PLF_2grFt_FH9_10[23] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[0]  (.D(\b13_PLF_2grFt_FH9_10[0] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(ttdo));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[6]  (.A(
        b8_FZFFLXYE[2]), .B(\b13_PLF_2grFt_FH9[7] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[6] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[11]  (.D(\b13_PLF_2grFt_FH9_10[11] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[11] ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[9]  (.A(
        b8_FZFFLXYE[5]), .B(\b13_PLF_2grFt_FH9[10] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[12]  (.D(\b13_PLF_2grFt_FH9_10[12] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[12] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[17]  (.D(\b13_PLF_2grFt_FH9_10[17] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[17] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[20]  (.D(\b13_PLF_2grFt_FH9_10[20] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[20] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[14]  (.D(\b13_PLF_2grFt_FH9_10[14] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[14] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[6]  (.D(\b13_PLF_2grFt_FH9_10[6] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[6] ));
    GND GND (.Y(GND_net_1));
    SLE \genblk1.b13_PLF_2grFt_FH9[21]  (.D(\b13_PLF_2grFt_FH9_10[21] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[21] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[17]  (.A(
        b12_PSyi_KyDbLbb[3]), .B(\b13_PLF_2grFt_FH9[18] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[17] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[20]  (.A(
        b12_PSyi_KyDbLbb[6]), .B(\b13_PLF_2grFt_FH9[21] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[20] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[22]  (.D(\b13_PLF_2grFt_FH9_10[22] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[22] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[18]  (.D(\b13_PLF_2grFt_FH9_10[18] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[18] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[21]  (.A(
        b12_PSyi_KyDbLbb[7]), .B(\b13_PLF_2grFt_FH9[22] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[21] ));
    CFG2 #( .INIT(4'h8) )  \genblk1.b13_PLF_2grFt_FH9_10[23]  (.A(
        IICE_comm2iice_4), .B(b12_PSyi_KyDbLbb[9]), .Y(
        \b13_PLF_2grFt_FH9_10[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[9]  (.D(\b13_PLF_2grFt_FH9_10[9] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[4]  (.D(\b13_PLF_2grFt_FH9_10[4] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[4] ));
    CFG4 #( .INIT(16'h8000) )  un1_b13_PLF_2grFt_FH923_i_a2 (.A(
        IICE_comm2iice_0), .B(un1_b13_PLF_2grFt_FH911_i_a2_0_1), .C(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .D(N_14_1), .Y(N_14));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[10]  (.A(
        b8_FZFFLXYE[6]), .B(\b13_PLF_2grFt_FH9[11] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[10] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[11]  (.A(
        b8_FZFFLXYE[7]), .B(\b13_PLF_2grFt_FH9[12] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[11] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[18]  (.A(
        b12_PSyi_KyDbLbb[4]), .B(\b13_PLF_2grFt_FH9[19] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[18] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[13]  (.A(
        b8_FZFFLXYE[9]), .B(\b13_PLF_2grFt_FH9[14] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[13] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[15]  (.D(\b13_PLF_2grFt_FH9_10[15] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[15] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[3]  (.D(\b13_PLF_2grFt_FH9_10[3] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[3] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[8]  (.A(
        b8_FZFFLXYE[4]), .B(\b13_PLF_2grFt_FH9[9] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[8] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[14]  (.A(
        b12_PSyi_KyDbLbb[0]), .B(\b13_PLF_2grFt_FH9[15] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[14] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[1]  (.D(\b13_PLF_2grFt_FH9_10[1] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[1] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[7]  (.D(\b13_PLF_2grFt_FH9_10[7] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[19]  (.D(\b13_PLF_2grFt_FH9_10[19] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[19] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[7]  (.A(
        b8_FZFFLXYE[3]), .B(\b13_PLF_2grFt_FH9[8] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[8]  (.D(\b13_PLF_2grFt_FH9_10[8] ), 
        .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[8] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[16]  (.A(
        b12_PSyi_KyDbLbb[2]), .B(\b13_PLF_2grFt_FH9[17] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[16] ));
    CFG3 #( .INIT(8'hAC) )  \genblk1.b13_PLF_2grFt_FH9_10[4]  (.A(
        b8_FZFFLXYE[0]), .B(\b13_PLF_2grFt_FH9[5] ), .C(
        IICE_comm2iice_4), .Y(\b13_PLF_2grFt_FH9_10[4] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[13]  (.D(\b13_PLF_2grFt_FH9_10[13] )
        , .CLK(IICE_comm2iice_6), .EN(N_14), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[13] ));
    
endmodule


module b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0(
       IICE_comm2iice_11,
       IICE_comm2iice_9,
       IICE_comm2iice_4,
       IICE_comm2iice_0,
       IICE_comm2iice_1,
       IICE_comm2iice_3,
       IICE_comm2iice_2,
       IICE_comm2iice_10,
       IICE_comm2iice_6,
       IICE_comm2iice_5,
       b4_ycsM,
       un1_b13_PLF_2grFt_FH911_i_a2_0_1,
       un1_b13_PLF_2grFt_FH911_i_a2_0_2,
       N_14_1
    );
input  IICE_comm2iice_11;
input  IICE_comm2iice_9;
input  IICE_comm2iice_4;
input  IICE_comm2iice_0;
input  IICE_comm2iice_1;
input  IICE_comm2iice_3;
input  IICE_comm2iice_2;
input  IICE_comm2iice_10;
input  IICE_comm2iice_6;
input  IICE_comm2iice_5;
output b4_ycsM;
output un1_b13_PLF_2grFt_FH911_i_a2_0_1;
output un1_b13_PLF_2grFt_FH911_i_a2_0_2;
output N_14_1;

    wire \b13_PLF_2grFt_FH9[24] , VCC_net_1, \b13_PLF_2grFt_FH9_5[24] , 
        N_13, GND_net_1, \b13_PLF_2grFt_FH9[25] , 
        \b13_PLF_2grFt_FH9_5[25] , \b13_PLF_2grFt_FH9[26] , 
        \b13_PLF_2grFt_FH9_5[26] , \b13_PLF_2grFt_FH9[27] , 
        \b13_PLF_2grFt_FH9_5[27] , \b13_PLF_2grFt_FH9[28] , 
        \b13_PLF_2grFt_FH9_5[28] , \b13_PLF_2grFt_FH9[29] , 
        \b13_PLF_2grFt_FH9_5[29] , \b13_PLF_2grFt_FH9[30] , 
        \b13_PLF_2grFt_FH9_5[30] , \b13_PLF_2grFt_FH9[31] , 
        \b13_PLF_2grFt_FH9[9] , \b13_PLF_2grFt_FH9_5[9] , 
        \b13_PLF_2grFt_FH9[10] , \b13_PLF_2grFt_FH9_5[10] , 
        \b13_PLF_2grFt_FH9[11] , \b13_PLF_2grFt_FH9_5[11] , 
        \b13_PLF_2grFt_FH9[12] , \b13_PLF_2grFt_FH9_5[12] , 
        \b13_PLF_2grFt_FH9[13] , \b13_PLF_2grFt_FH9_5[13] , 
        \b13_PLF_2grFt_FH9[14] , \b13_PLF_2grFt_FH9_5[14] , 
        \b13_PLF_2grFt_FH9[15] , \b13_PLF_2grFt_FH9_5[15] , 
        \b13_PLF_2grFt_FH9[16] , \b13_PLF_2grFt_FH9_5[16] , 
        \b13_PLF_2grFt_FH9[17] , \b13_PLF_2grFt_FH9_5[17] , 
        \b13_PLF_2grFt_FH9[18] , \b13_PLF_2grFt_FH9_5[18] , 
        \b13_PLF_2grFt_FH9[19] , \b13_PLF_2grFt_FH9_5[19] , 
        \b13_PLF_2grFt_FH9[20] , \b13_PLF_2grFt_FH9_5[20] , 
        \b13_PLF_2grFt_FH9[21] , \b13_PLF_2grFt_FH9_5[21] , 
        \b13_PLF_2grFt_FH9[22] , \b13_PLF_2grFt_FH9_5[22] , 
        \b13_PLF_2grFt_FH9[23] , \b13_PLF_2grFt_FH9_5[23] , 
        \b13_PLF_2grFt_FH9_5[0] , \b13_PLF_2grFt_FH9[1] , 
        \b13_PLF_2grFt_FH9_5[1] , \b13_PLF_2grFt_FH9[2] , 
        \b13_PLF_2grFt_FH9_5[2] , \b13_PLF_2grFt_FH9[3] , 
        \b13_PLF_2grFt_FH9_5[3] , \b13_PLF_2grFt_FH9[4] , 
        \b13_PLF_2grFt_FH9_5[4] , \b13_PLF_2grFt_FH9[5] , 
        \b13_PLF_2grFt_FH9_5[5] , \b13_PLF_2grFt_FH9[6] , 
        \b13_PLF_2grFt_FH9_5[6] , \b13_PLF_2grFt_FH9[7] , 
        \b13_PLF_2grFt_FH9_5[7] , \b13_PLF_2grFt_FH9[8] , 
        \b13_PLF_2grFt_FH9_5[8] ;
    
    SLE \genblk1.b13_PLF_2grFt_FH9[2]  (.D(\b13_PLF_2grFt_FH9_5[2] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[2] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[22]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[23] ), .Y(
        \b13_PLF_2grFt_FH9_5[22] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[26]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[27] ), .Y(
        \b13_PLF_2grFt_FH9_5[26] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[5]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[6] ), .Y(
        \b13_PLF_2grFt_FH9_5[5] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[5]  (.D(\b13_PLF_2grFt_FH9_5[5] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[5] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[16]  (.D(\b13_PLF_2grFt_FH9_5[16] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[16] ));
    CFG3 #( .INIT(8'h20) )  un1_b13_PLF_2grFt_FH911_i_a2_0_2_inst_1 (
        .A(IICE_comm2iice_1), .B(IICE_comm2iice_3), .C(
        IICE_comm2iice_2), .Y(un1_b13_PLF_2grFt_FH911_i_a2_0_2));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[3]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[4] ), .Y(
        \b13_PLF_2grFt_FH9_5[3] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[10]  (.D(\b13_PLF_2grFt_FH9_5[10] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[10] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[25]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[26] ), .Y(
        \b13_PLF_2grFt_FH9_5[25] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[23]  (.D(\b13_PLF_2grFt_FH9_5[23] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[0]  (.D(\b13_PLF_2grFt_FH9_5[0] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b4_ycsM));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[30]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[31] ), .Y(
        \b13_PLF_2grFt_FH9_5[30] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[20]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[21] ), .Y(
        \b13_PLF_2grFt_FH9_5[20] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[11]  (.D(\b13_PLF_2grFt_FH9_5[11] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[11] ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[21]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[22] ), .Y(
        \b13_PLF_2grFt_FH9_5[21] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[18]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[19] ), .Y(
        \b13_PLF_2grFt_FH9_5[18] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[1]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[2] ), .Y(
        \b13_PLF_2grFt_FH9_5[1] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[12]  (.D(\b13_PLF_2grFt_FH9_5[12] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[12] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[17]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[18] ), .Y(
        \b13_PLF_2grFt_FH9_5[17] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[4]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[5] ), .Y(
        \b13_PLF_2grFt_FH9_5[4] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[17]  (.D(\b13_PLF_2grFt_FH9_5[17] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[17] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[26]  (.D(\b13_PLF_2grFt_FH9_5[26] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[26] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[20]  (.D(\b13_PLF_2grFt_FH9_5[20] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[20] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[24]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[25] ), .Y(
        \b13_PLF_2grFt_FH9_5[24] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[13]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[14] ), .Y(
        \b13_PLF_2grFt_FH9_5[13] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[14]  (.D(\b13_PLF_2grFt_FH9_5[14] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[14] ));
    CFG3 #( .INIT(8'hE0) )  un1_b13_PLF_2grFt_FH911_i_a2_1_0 (.A(
        IICE_comm2iice_9), .B(IICE_comm2iice_10), .C(IICE_comm2iice_6), 
        .Y(N_14_1));
    CFG2 #( .INIT(4'h4) )  un1_b13_PLF_2grFt_FH911_i_a2_0_1_inst_1 (.A(
        IICE_comm2iice_4), .B(IICE_comm2iice_0), .Y(
        un1_b13_PLF_2grFt_FH911_i_a2_0_1));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[29]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[30] ), .Y(
        \b13_PLF_2grFt_FH9_5[29] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[6]  (.D(\b13_PLF_2grFt_FH9_5[6] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[6] ));
    GND GND (.Y(GND_net_1));
    SLE \genblk1.b13_PLF_2grFt_FH9[21]  (.D(\b13_PLF_2grFt_FH9_5[21] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[21] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[0]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[1] ), .Y(
        \b13_PLF_2grFt_FH9_5[0] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[22]  (.D(\b13_PLF_2grFt_FH9_5[22] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[22] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[18]  (.D(\b13_PLF_2grFt_FH9_5[18] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[18] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[12]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[13] ), .Y(
        \b13_PLF_2grFt_FH9_5[12] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[16]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[17] ), .Y(
        \b13_PLF_2grFt_FH9_5[16] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[9]  (.D(\b13_PLF_2grFt_FH9_5[9] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[4]  (.D(\b13_PLF_2grFt_FH9_5[4] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[4] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[27]  (.D(\b13_PLF_2grFt_FH9_5[27] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[27] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[30]  (.D(\b13_PLF_2grFt_FH9_5[30] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[30] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[8]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[9] ), .Y(
        \b13_PLF_2grFt_FH9_5[8] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[24]  (.D(\b13_PLF_2grFt_FH9_5[24] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[24] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[15]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[16] ), .Y(
        \b13_PLF_2grFt_FH9_5[15] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[15]  (.D(\b13_PLF_2grFt_FH9_5[15] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[15] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[10]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[11] ), .Y(
        \b13_PLF_2grFt_FH9_5[10] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[3]  (.D(\b13_PLF_2grFt_FH9_5[3] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[3] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[31]  (.D(IICE_comm2iice_9), .CLK(
        IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b13_PLF_2grFt_FH9[31] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[9]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[10] ), .Y(
        \b13_PLF_2grFt_FH9_5[9] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[1]  (.D(\b13_PLF_2grFt_FH9_5[1] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[1] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[11]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[12] ), .Y(
        \b13_PLF_2grFt_FH9_5[11] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[7]  (.D(\b13_PLF_2grFt_FH9_5[7] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[19]  (.D(\b13_PLF_2grFt_FH9_5[19] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[19] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[6]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[7] ), .Y(
        \b13_PLF_2grFt_FH9_5[6] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[7]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[8] ), .Y(
        \b13_PLF_2grFt_FH9_5[7] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[28]  (.D(\b13_PLF_2grFt_FH9_5[28] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[28] ));
    CFG2 #( .INIT(4'h4) )  \genblk1.b13_PLF_2grFt_FH9_5[28]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[29] ), .Y(
        \b13_PLF_2grFt_FH9_5[28] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[8]  (.D(\b13_PLF_2grFt_FH9_5[8] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[8] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[27]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[28] ), .Y(
        \b13_PLF_2grFt_FH9_5[27] ));
    CFG4 #( .INIT(16'h4000) )  un1_b13_PLF_2grFt_FH911_i_a2 (.A(
        IICE_comm2iice_5), .B(un1_b13_PLF_2grFt_FH911_i_a2_0_1), .C(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .D(N_14_1), .Y(N_13));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[14]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[15] ), .Y(
        \b13_PLF_2grFt_FH9_5[14] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[2]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[3] ), .Y(
        \b13_PLF_2grFt_FH9_5[2] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[25]  (.D(\b13_PLF_2grFt_FH9_5[25] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[25] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[19]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[20] ), .Y(
        \b13_PLF_2grFt_FH9_5[19] ));
    CFG2 #( .INIT(4'hE) )  \genblk1.b13_PLF_2grFt_FH9_5[23]  (.A(
        IICE_comm2iice_9), .B(\b13_PLF_2grFt_FH9[24] ), .Y(
        \b13_PLF_2grFt_FH9_5[23] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[29]  (.D(\b13_PLF_2grFt_FH9_5[29] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[29] ));
    SLE \genblk1.b13_PLF_2grFt_FH9[13]  (.D(\b13_PLF_2grFt_FH9_5[13] ), 
        .CLK(IICE_comm2iice_11), .EN(N_13), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b13_PLF_2grFt_FH9[13] ));
    
endmodule


module b11_SoWyP0zEFKY_161s_0s_6s_0s_2s_2s_0s_0s_2s_0s_x_0(
       b11_OFWNT9L_8tZ,
       mdiclink_reg,
       b13_nAzGfFM_sLsv3,
       BW_clk_c,
       b8_SoWGfWYY,
       b4_2o_z,
       b13_oRB_MqCD2_EdR_RNI9OIA,
       N_44
    );
output [154:0] b11_OFWNT9L_8tZ;
input  [154:0] mdiclink_reg;
input  [1:1] b13_nAzGfFM_sLsv3;
input  BW_clk_c;
input  b8_SoWGfWYY;
output b4_2o_z;
output b13_oRB_MqCD2_EdR_RNI9OIA;
input  N_44;

    wire VCC_net_1, GND_net_1, b13_oRB_MqCD2_EdR;
    
    SLE \genblk2.b5_oRB_C[72]  (.D(mdiclink_reg[82]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[72]));
    SLE \genblk2.b5_oRB_C[61]  (.D(mdiclink_reg[93]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[61]));
    SLE \genblk2.b5_oRB_C[131]  (.D(mdiclink_reg[23]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[131]));
    SLE \genblk2.b5_oRB_C[82]  (.D(mdiclink_reg[72]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[82]));
    SLE \genblk2.b5_oRB_C[122]  (.D(mdiclink_reg[32]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[122]));
    SLE \genblk2.b5_oRB_C[17]  (.D(mdiclink_reg[137]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[17]));
    SLE \genblk2.b5_oRB_C[18]  (.D(mdiclink_reg[136]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[18]));
    SLE \genblk2.b5_oRB_C[66]  (.D(mdiclink_reg[88]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[66]));
    SLE \genblk2.b5_oRB_C[137]  (.D(mdiclink_reg[17]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[137]));
    SLE \genblk2.b5_oRB_C[105]  (.D(mdiclink_reg[49]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[105]));
    SLE \genblk2.b5_oRB_C[121]  (.D(mdiclink_reg[33]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[121]));
    SLE \genblk2.b5_oRB_C[20]  (.D(mdiclink_reg[134]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[20]));
    SLE \genblk2.b5_oRB_C[43]  (.D(mdiclink_reg[111]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[43]));
    SLE \genblk2.b5_oRB_C[93]  (.D(mdiclink_reg[61]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[93]));
    SLE \genblk2.b5_oRB_C[11]  (.D(mdiclink_reg[143]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[11]));
    SLE \genblk2.b5_oRB_C[127]  (.D(mdiclink_reg[27]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[127]));
    SLE \genblk2.b5_oRB_C[30]  (.D(mdiclink_reg[124]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[30]));
    SLE \genblk2.b5_oRB_C[16]  (.D(mdiclink_reg[138]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[16]));
    SLE \genblk2.b5_oRB_C[45]  (.D(mdiclink_reg[109]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[45]));
    SLE \genblk2.b5_oRB_C[95]  (.D(mdiclink_reg[59]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[95]));
    SLE \genblk2.b5_oRB_C[70]  (.D(mdiclink_reg[84]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[70]));
    SLE \genblk2.b5_oRB_C[5]  (.D(mdiclink_reg[149]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[5]));
    SLE \genblk2.b5_oRB_C[80]  (.D(mdiclink_reg[74]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[80]));
    SLE \genblk2.b5_oRB_C[0]  (.D(mdiclink_reg[154]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[0]));
    SLE \genblk2.b5_oRB_C[104]  (.D(mdiclink_reg[50]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[104]));
    SLE \genblk2.b5_oRB_C[57]  (.D(mdiclink_reg[97]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[57]));
    SLE \genblk2.b5_oRB_C[58]  (.D(mdiclink_reg[96]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[58]));
    SLE \genblk2.b5_oRB_C[63]  (.D(mdiclink_reg[91]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[63]));
    SLE \genblk2.b5_oRB_C[106]  (.D(mdiclink_reg[48]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[106]));
    SLE \genblk2.b5_oRB_C[65]  (.D(mdiclink_reg[89]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[65]));
    GND GND (.Y(GND_net_1));
    SLE \genblk2.b5_oRB_C[51]  (.D(mdiclink_reg[103]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[51]));
    SLE \genblk2.b5_oRB_C[115]  (.D(mdiclink_reg[39]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[115]));
    SLE \genblk2.b5_oRB_C[13]  (.D(mdiclink_reg[141]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[13]));
    SLE \genblk2.b5_oRB_C[56]  (.D(mdiclink_reg[98]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[56]));
    SLE \genblk2.b5_oRB_C[44]  (.D(mdiclink_reg[110]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[44]));
    SLE \genblk2.b5_oRB_C[94]  (.D(mdiclink_reg[60]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[94]));
    SLE \genblk2.b5_oRB_C[15]  (.D(mdiclink_reg[139]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[15]));
    CFG2 #( .INIT(4'hE) )  \genblk2.b13_oRB_MqCD2_EdR_RNI9OIA  (.A(
        b8_SoWGfWYY), .B(b4_2o_z), .Y(b13_oRB_MqCD2_EdR_RNI9OIA));
    SLE \genblk2.b5_oRB_C[3]  (.D(mdiclink_reg[151]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[3]));
    SLE \genblk2.b5_oRB_C[114]  (.D(mdiclink_reg[40]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[114]));
    SLE \genblk2.b5_oRB_C[108]  (.D(mdiclink_reg[46]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[108]));
    SLE \genblk2.b5_oRB_C[154]  (.D(mdiclink_reg[0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[154]));
    SLE \genblk2.b5_oRB_C[53]  (.D(mdiclink_reg[101]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[53]));
    SLE \genblk2.b5_oRB_C[64]  (.D(mdiclink_reg[90]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[64]));
    SLE \genblk2.b5_oRB_C[116]  (.D(mdiclink_reg[38]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[116]));
    SLE \genblk2.b5_oRB_C[49]  (.D(mdiclink_reg[105]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[49]));
    SLE \genblk2.b5_oRB_C[99]  (.D(mdiclink_reg[55]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[99]));
    VCC VCC (.Y(VCC_net_1));
    SLE \genblk2.b5_oRB_C[100]  (.D(mdiclink_reg[54]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[100]));
    SLE \genblk2.b5_oRB_C[103]  (.D(mdiclink_reg[51]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[103]));
    SLE \genblk2.b5_oRB_C[145]  (.D(mdiclink_reg[9]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[145]));
    SLE \genblk2.b5_oRB_C[55]  (.D(mdiclink_reg[99]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[55]));
    SLE \genblk2.b5_oRB_C[27]  (.D(mdiclink_reg[127]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[27]));
    SLE \genblk2.b5_oRB_C[28]  (.D(mdiclink_reg[126]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[28]));
    SLE \genblk2.b5_oRB_C[14]  (.D(mdiclink_reg[140]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[14]));
    SLE \genblk2.b5_oRB_C[37]  (.D(mdiclink_reg[117]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[37]));
    SLE \genblk2.b5_oRB_C[38]  (.D(mdiclink_reg[116]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[38]));
    SLE \genblk2.b5_oRB_C[69]  (.D(mdiclink_reg[85]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[69]));
    SLE \genblk2.b5_oRB_C[109]  (.D(mdiclink_reg[45]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[109]));
    SLE \genblk2.b5_oRB_C[1]  (.D(mdiclink_reg[153]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[1]));
    SLE \genblk2.b5_oRB_C[21]  (.D(mdiclink_reg[133]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[21]));
    SLE \genblk2.b5_oRB_C[77]  (.D(mdiclink_reg[77]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[77]));
    SLE \genblk2.b5_oRB_C[144]  (.D(mdiclink_reg[10]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[144]));
    SLE \genblk2.b5_oRB_C[78]  (.D(mdiclink_reg[76]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[78]));
    SLE \genblk2.b5_oRB_C[87]  (.D(mdiclink_reg[67]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[87]));
    SLE \genblk2.b5_oRB_C[88]  (.D(mdiclink_reg[66]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[88]));
    SLE \genblk2.b5_oRB_C[42]  (.D(mdiclink_reg[112]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[42]));
    SLE \genblk2.b5_oRB_C[92]  (.D(mdiclink_reg[62]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[92]));
    SLE \genblk2.b5_oRB_C[118]  (.D(mdiclink_reg[36]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[118]));
    SLE \genblk2.b5_oRB_C[26]  (.D(mdiclink_reg[128]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[26]));
    SLE \genblk2.b5_oRB_C[31]  (.D(mdiclink_reg[123]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[31]));
    SLE \genblk2.b5_oRB_C[36]  (.D(mdiclink_reg[118]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[36]));
    SLE \genblk2.b5_oRB_C[146]  (.D(mdiclink_reg[8]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[146]));
    SLE \genblk2.b5_oRB_C[19]  (.D(mdiclink_reg[135]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[19]));
    SLE \genblk2.b5_oRB_C[9]  (.D(mdiclink_reg[145]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[9]));
    SLE \genblk2.b5_oRB_C[71]  (.D(mdiclink_reg[83]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[71]));
    SLE \genblk2.b5_oRB_C[102]  (.D(mdiclink_reg[52]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[102]));
    SLE \genblk2.b5_oRB_C[54]  (.D(mdiclink_reg[100]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[54]));
    SLE \genblk2.b5_oRB_C[81]  (.D(mdiclink_reg[73]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[81]));
    SLE \genblk2.b5_oRB_C[110]  (.D(mdiclink_reg[44]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[110]));
    SLE \genblk2.b5_oRB_C[113]  (.D(mdiclink_reg[41]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[113]));
    SLE \genblk2.b5_oRB_C[76]  (.D(mdiclink_reg[78]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[76]));
    SLE \genblk2.b5_oRB_C[86]  (.D(mdiclink_reg[68]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[86]));
    SLE \genblk2.b5_oRB_C[150]  (.D(mdiclink_reg[4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[150]));
    SLE \genblk2.b5_oRB_C[153]  (.D(mdiclink_reg[1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[153]));
    SLE \genblk2.b5_oRB_C[101]  (.D(mdiclink_reg[53]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[101]));
    SLE \genblk2.b5_oRB_C[62]  (.D(mdiclink_reg[92]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[62]));
    SLE \genblk2.b5_oRB_C[135]  (.D(mdiclink_reg[19]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[135]));
    SLE \genblk2.b13_oRB_MqCD2_EdR  (.D(b13_oRB_MqCD2_EdR), .CLK(
        BW_clk_c), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(b4_2o_z));
    SLE \genblk2.b5_oRB_C[40]  (.D(mdiclink_reg[114]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[40]));
    SLE \genblk2.b5_oRB_C[107]  (.D(mdiclink_reg[47]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[107]));
    SLE \genblk2.b5_oRB_C[90]  (.D(mdiclink_reg[64]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[90]));
    SLE \genblk2.b5_oRB_C[23]  (.D(mdiclink_reg[131]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[23]));
    SLE \genblk2.b5_oRB_C[125]  (.D(mdiclink_reg[29]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[125]));
    SLE \genblk2.b5_oRB_C[119]  (.D(mdiclink_reg[35]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[119]));
    SLE \genblk2.b5_oRB_C[33]  (.D(mdiclink_reg[121]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[33]));
    SLE \genblk2.b5_oRB_C[59]  (.D(mdiclink_reg[95]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[59]));
    SLE \genblk2.b5_oRB_C[12]  (.D(mdiclink_reg[142]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[12]));
    SLE \genblk2.b5_oRB_C[7]  (.D(mdiclink_reg[147]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[7]));
    SLE \genblk2.b5_oRB_C[25]  (.D(mdiclink_reg[129]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[25]));
    SLE \genblk2.b5_oRB_C[148]  (.D(mdiclink_reg[6]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[148]));
    SLE \genblk2.b5_oRB_C[134]  (.D(mdiclink_reg[20]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[134]));
    SLE \genblk2.b5_oRB_C[73]  (.D(mdiclink_reg[81]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[73]));
    SLE \genblk2.b5_oRB_C[83]  (.D(mdiclink_reg[71]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[83]));
    SLE \genblk2.b5_oRB_C[35]  (.D(mdiclink_reg[119]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[35]));
    SLE \genblk2.b5_oRB_C[60]  (.D(mdiclink_reg[94]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[60]));
    SLE \genblk2.b5_oRB_C[112]  (.D(mdiclink_reg[42]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[112]));
    SLE \genblk2.b5_oRB_C[140]  (.D(mdiclink_reg[14]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[140]));
    SLE \genblk2.b5_oRB_C[143]  (.D(mdiclink_reg[11]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[143]));
    SLE \genblk2.b5_oRB_C[124]  (.D(mdiclink_reg[30]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[124]));
    SLE \genblk2.b5_oRB_C[75]  (.D(mdiclink_reg[79]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[75]));
    SLE \genblk2.b5_oRB_C[136]  (.D(mdiclink_reg[18]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[136]));
    SLE \genblk2.b5_oRB_C[85]  (.D(mdiclink_reg[69]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[85]));
    SLE \genblk2.b5_oRB_C[152]  (.D(mdiclink_reg[2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[152]));
    SLE \genblk2.b5_oRB_C[111]  (.D(mdiclink_reg[43]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[111]));
    SLE \genblk2.b5_oRB_C[8]  (.D(mdiclink_reg[146]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[8]));
    SLE \genblk2.b5_oRB_C[2]  (.D(mdiclink_reg[152]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[2]));
    SLE \genblk2.b5_oRB_C[126]  (.D(mdiclink_reg[28]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[126]));
    SLE \genblk2.b5_oRB_C[10]  (.D(mdiclink_reg[144]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[10]));
    SLE \genblk2.b5_oRB_C[52]  (.D(mdiclink_reg[102]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[52]));
    SLE \genblk2.b5_oRB_C[151]  (.D(mdiclink_reg[3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[151]));
    SLE \genblk2.b5_oRB_C[117]  (.D(mdiclink_reg[37]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[117]));
    SLE \genblk2.b5_oRB_C[149]  (.D(mdiclink_reg[5]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[149]));
    SLE \genblk2.b5_oRB_C[24]  (.D(mdiclink_reg[130]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[24]));
    CFG2 #( .INIT(4'hE) )  \genblk2.b13_oRB_MqCD2_EdR_s  (.A(N_44), .B(
        b13_nAzGfFM_sLsv3[1]), .Y(b13_oRB_MqCD2_EdR));
    SLE \genblk2.b5_oRB_C[34]  (.D(mdiclink_reg[120]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[34]));
    SLE \genblk2.b5_oRB_C[4]  (.D(mdiclink_reg[150]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[4]));
    SLE \genblk2.b5_oRB_C[138]  (.D(mdiclink_reg[16]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[138]));
    SLE \genblk2.b5_oRB_C[142]  (.D(mdiclink_reg[12]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[142]));
    SLE \genblk2.b5_oRB_C[74]  (.D(mdiclink_reg[80]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[74]));
    SLE \genblk2.b5_oRB_C[84]  (.D(mdiclink_reg[70]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[84]));
    SLE \genblk2.b5_oRB_C[50]  (.D(mdiclink_reg[104]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[50]));
    SLE \genblk2.b5_oRB_C[128]  (.D(mdiclink_reg[26]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[128]));
    SLE \genblk2.b5_oRB_C[130]  (.D(mdiclink_reg[24]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[130]));
    SLE \genblk2.b5_oRB_C[141]  (.D(mdiclink_reg[13]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[141]));
    SLE \genblk2.b5_oRB_C[133]  (.D(mdiclink_reg[21]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[133]));
    SLE \genblk2.b5_oRB_C[29]  (.D(mdiclink_reg[125]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[29]));
    SLE \genblk2.b5_oRB_C[147]  (.D(mdiclink_reg[7]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[147]));
    SLE \genblk2.b5_oRB_C[39]  (.D(mdiclink_reg[115]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[39]));
    SLE \genblk2.b5_oRB_C[120]  (.D(mdiclink_reg[34]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[120]));
    SLE \genblk2.b5_oRB_C[123]  (.D(mdiclink_reg[31]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[123]));
    SLE \genblk2.b5_oRB_C[47]  (.D(mdiclink_reg[107]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[47]));
    SLE \genblk2.b5_oRB_C[97]  (.D(mdiclink_reg[57]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[97]));
    SLE \genblk2.b5_oRB_C[48]  (.D(mdiclink_reg[106]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[48]));
    SLE \genblk2.b5_oRB_C[98]  (.D(mdiclink_reg[56]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[98]));
    SLE \genblk2.b5_oRB_C[79]  (.D(mdiclink_reg[75]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[79]));
    SLE \genblk2.b5_oRB_C[89]  (.D(mdiclink_reg[65]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[89]));
    SLE \genblk2.b5_oRB_C[139]  (.D(mdiclink_reg[15]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[139]));
    SLE \genblk2.b5_oRB_C[6]  (.D(mdiclink_reg[148]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[6]));
    SLE \genblk2.b5_oRB_C[41]  (.D(mdiclink_reg[113]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[41]));
    SLE \genblk2.b5_oRB_C[91]  (.D(mdiclink_reg[63]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[91]));
    SLE \genblk2.b5_oRB_C[129]  (.D(mdiclink_reg[25]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[129]));
    SLE \genblk2.b5_oRB_C[22]  (.D(mdiclink_reg[132]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[22]));
    SLE \genblk2.b5_oRB_C[46]  (.D(mdiclink_reg[108]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[46]));
    SLE \genblk2.b5_oRB_C[96]  (.D(mdiclink_reg[58]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[96]));
    SLE \genblk2.b5_oRB_C[67]  (.D(mdiclink_reg[87]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[67]));
    SLE \genblk2.b5_oRB_C[68]  (.D(mdiclink_reg[86]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[68]));
    SLE \genblk2.b5_oRB_C[32]  (.D(mdiclink_reg[122]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[32]));
    SLE \genblk2.b5_oRB_C[132]  (.D(mdiclink_reg[22]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b11_OFWNT9L_8tZ[132]));
    
endmodule


module b11_OFWNT9s_8tZ_Z2_x(
       b11_OFWNT9L_8tZ,
       mdiclink_reg,
       b13_nAzGfFM_sLsv3,
       IICE_comm2iice_11,
       IICE_comm2iice_0,
       IICE_comm2iice_4,
       IICE_comm2iice_10,
       IICE_comm2iice_5,
       IICE_comm2iice_9,
       IICE_comm2iice_1,
       IICE_comm2iice_3,
       IICE_comm2iice_2,
       IICE_comm2iice_6,
       BW_clk_c,
       b11_PSyil9s_FMZ,
       b8_SoWGfWYY_i,
       b8_SoWGfWYY,
       b7_yYh03wy,
       b10_OFWNT9khFt,
       b9_OFWNT9Mxf,
       N_44
    );
output [154:0] b11_OFWNT9L_8tZ;
input  [154:0] mdiclink_reg;
input  [1:1] b13_nAzGfFM_sLsv3;
input  IICE_comm2iice_11;
input  IICE_comm2iice_0;
input  IICE_comm2iice_4;
input  IICE_comm2iice_10;
input  IICE_comm2iice_5;
input  IICE_comm2iice_9;
input  IICE_comm2iice_1;
input  IICE_comm2iice_3;
input  IICE_comm2iice_2;
input  IICE_comm2iice_6;
input  BW_clk_c;
input  b11_PSyil9s_FMZ;
input  b8_SoWGfWYY_i;
input  b8_SoWGfWYY;
output b7_yYh03wy;
input  b10_OFWNT9khFt;
output b9_OFWNT9Mxf;
input  N_44;

    wire \b12_PSyi_KyDbLbb[1]_net_1 , VCC_net_1, 
        \b12_2_St6KCa_jHv[1]_net_1 , b12_PSyi_KyDbLbb_0_sqmuxa_net_1, 
        GND_net_1, \b12_PSyi_KyDbLbb[2]_net_1 , 
        \b12_2_St6KCa_jHv[2]_net_1 , \b12_PSyi_KyDbLbb[3]_net_1 , 
        \b12_2_St6KCa_jHv[3]_net_1 , \b12_PSyi_KyDbLbb[4]_net_1 , 
        \b12_2_St6KCa_jHv[4]_net_1 , \b12_PSyi_KyDbLbb[5]_net_1 , 
        \b12_2_St6KCa_jHv[5]_net_1 , \b12_PSyi_KyDbLbb[6]_net_1 , 
        \b12_2_St6KCa_jHv[6]_net_1 , \b12_PSyi_KyDbLbb[7]_net_1 , 
        \b12_2_St6KCa_jHv[7]_net_1 , \b12_PSyi_KyDbLbb[8]_net_1 , 
        \b12_2_St6KCa_jHv[8]_net_1 , \b12_PSyi_KyDbLbb[9]_net_1 , 
        \b12_2_St6KCa_jHv[9]_net_1 , \b12_PSyi_KyDbLbb[0]_net_1 , 
        \b12_2_St6KCa_jHv[0]_net_1 , b9_PSyil9s_2_net_1, b8_nYJ_TqLY, 
        \b7_nYJ_BFM[160] , \b7_nYJ_BFM_or[10] , \b7_nYJ_BFM[146] , 
        \b7_nYJ_BFM[145] , \b7_nYJ_BFM[147] , \b7_nYJ_BFM[148] , 
        \b7_nYJ_BFM[149] , \b7_nYJ_BFM[150] , \b7_nYJ_BFM[151] , 
        \b7_nYJ_BFM[152] , \b7_nYJ_BFM[153] , \b7_nYJ_BFM[154] , 
        \b7_nYJ_BFM[155] , \b7_nYJ_BFM[156] , \b7_nYJ_BFM[157] , 
        \b7_nYJ_BFM[158] , \b7_nYJ_BFM[159] , \b7_nYJ_BFM[131] , 
        \b7_nYJ_BFM[130] , \b7_nYJ_BFM[132] , \b7_nYJ_BFM[133] , 
        \b7_nYJ_BFM[134] , \b7_nYJ_BFM[135] , \b7_nYJ_BFM[136] , 
        \b7_nYJ_BFM[137] , \b7_nYJ_BFM[138] , \b7_nYJ_BFM[139] , 
        \b7_nYJ_BFM[140] , \b7_nYJ_BFM[141] , \b7_nYJ_BFM[142] , 
        \b7_nYJ_BFM[143] , \b7_nYJ_BFM[144] , \b7_nYJ_BFM[116] , 
        \b7_nYJ_BFM[115] , \b7_nYJ_BFM[117] , \b7_nYJ_BFM[118] , 
        \b7_nYJ_BFM[119] , \b7_nYJ_BFM[120] , \b7_nYJ_BFM[121] , 
        \b7_nYJ_BFM[122] , \b7_nYJ_BFM[123] , \b7_nYJ_BFM[124] , 
        \b7_nYJ_BFM[125] , \b7_nYJ_BFM[126] , \b7_nYJ_BFM[127] , 
        \b7_nYJ_BFM[128] , \b7_nYJ_BFM[129] , \b7_nYJ_BFM[101] , 
        \b7_nYJ_BFM[100] , \b7_nYJ_BFM[102] , \b7_nYJ_BFM[103] , 
        \b7_nYJ_BFM[104] , \b7_nYJ_BFM[105] , \b7_nYJ_BFM[106] , 
        \b7_nYJ_BFM[107] , \b7_nYJ_BFM[108] , \b7_nYJ_BFM[109] , 
        \b7_nYJ_BFM[110] , \b7_nYJ_BFM[111] , \b7_nYJ_BFM[112] , 
        \b7_nYJ_BFM[113] , \b7_nYJ_BFM[114] , \b7_nYJ_BFM[86] , 
        \b7_nYJ_BFM[85] , \b7_nYJ_BFM[87] , \b7_nYJ_BFM[88] , 
        \b7_nYJ_BFM[89] , \b7_nYJ_BFM[90] , \b7_nYJ_BFM[91] , 
        \b7_nYJ_BFM[92] , \b7_nYJ_BFM[93] , \b7_nYJ_BFM[94] , 
        \b7_nYJ_BFM[95] , \b7_nYJ_BFM[96] , \b7_nYJ_BFM[97] , 
        \b7_nYJ_BFM[98] , \b7_nYJ_BFM[99] , \b7_nYJ_BFM[71] , 
        \b7_nYJ_BFM[70] , \b7_nYJ_BFM[72] , \b7_nYJ_BFM[73] , 
        \b7_nYJ_BFM[74] , \b7_nYJ_BFM[75] , \b7_nYJ_BFM[76] , 
        \b7_nYJ_BFM[77] , \b7_nYJ_BFM[78] , \b7_nYJ_BFM[79] , 
        \b7_nYJ_BFM[80] , \b7_nYJ_BFM[81] , \b7_nYJ_BFM[82] , 
        \b7_nYJ_BFM[83] , \b7_nYJ_BFM[84] , \b7_nYJ_BFM[56] , 
        \b7_nYJ_BFM[55] , \b7_nYJ_BFM[57] , \b7_nYJ_BFM[58] , 
        \b7_nYJ_BFM[59] , \b7_nYJ_BFM[60] , \b7_nYJ_BFM[61] , 
        \b7_nYJ_BFM[62] , \b7_nYJ_BFM[63] , \b7_nYJ_BFM[64] , 
        \b7_nYJ_BFM[65] , \b7_nYJ_BFM[66] , \b7_nYJ_BFM[67] , 
        \b7_nYJ_BFM[68] , \b7_nYJ_BFM[69] , \b7_nYJ_BFM[41] , 
        \b7_nYJ_BFM[40] , \b7_nYJ_BFM[42] , \b7_nYJ_BFM[43] , 
        \b7_nYJ_BFM[44] , \b7_nYJ_BFM[45] , \b7_nYJ_BFM[46] , 
        \b7_nYJ_BFM[47] , \b7_nYJ_BFM[48] , \b7_nYJ_BFM[49] , 
        \b7_nYJ_BFM[50] , \b7_nYJ_BFM[51] , \b7_nYJ_BFM[52] , 
        \b7_nYJ_BFM[53] , \b7_nYJ_BFM[54] , \b7_nYJ_BFM[26] , 
        \b7_nYJ_BFM[25] , \b7_nYJ_BFM[27] , \b7_nYJ_BFM[28] , 
        \b7_nYJ_BFM[29] , \b7_nYJ_BFM[30] , \b7_nYJ_BFM[31] , 
        \b7_nYJ_BFM[32] , \b7_nYJ_BFM[33] , \b7_nYJ_BFM[34] , 
        \b7_nYJ_BFM[35] , \b7_nYJ_BFM[36] , \b7_nYJ_BFM[37] , 
        \b7_nYJ_BFM[38] , \b7_nYJ_BFM[39] , \b7_nYJ_BFM[11] , 
        \b7_nYJ_BFM[10] , \b7_nYJ_BFM[12] , \b7_nYJ_BFM[13] , 
        \b7_nYJ_BFM[14] , \b7_nYJ_BFM[15] , \b7_nYJ_BFM[16] , 
        \b7_nYJ_BFM[17] , \b7_nYJ_BFM[18] , \b7_nYJ_BFM[19] , 
        \b7_nYJ_BFM[20] , \b7_nYJ_BFM[21] , \b7_nYJ_BFM[22] , 
        \b7_nYJ_BFM[23] , \b7_nYJ_BFM[24] , \b8_FZFFLXYE[6]_net_1 , 
        b13_oRB_MqCD2_EdR_RNI9OIA, \b8_FZFFLXYE[7]_net_1 , 
        \b8_FZFFLXYE[8]_net_1 , \b8_FZFFLXYE[9]_net_1 , 
        \b7_nYJ_BFM[0] , \b7_nYJ_BFM[1] , \b7_nYJ_BFM[2] , 
        \b7_nYJ_BFM[3] , \b7_nYJ_BFM[4] , \b7_nYJ_BFM[5] , 
        \b7_nYJ_BFM[6] , \b7_nYJ_BFM[7] , \b7_nYJ_BFM[8] , 
        \b7_nYJ_BFM[9] , N_406_a2_1_net_1, \b8_FZFFLXYE[0]_net_1 , 
        \b8_FZFFLXYE[1]_net_1 , \b8_FZFFLXYE[2]_net_1 , 
        \b8_FZFFLXYE[3]_net_1 , \b8_FZFFLXYE[4]_net_1 , 
        \b8_FZFFLXYE[5]_net_1 , b8_jAA_KlCO_net_1, 
        b8_jAA_KlCO_RNO_net_1, b8_jAA_KlCO_0_sqmuxa_net_1, 
        \b9_v_mzCDYXs[4] , b9_v_mzCDYXs_8, \b9_v_mzCDYXs[5] , 
        b9_v_mzCDYXs_7, \b9_v_mzCDYXs[6] , b9_v_mzCDYXs_6, 
        \b9_v_mzCDYXs[7] , b9_v_mzCDYXs_5, \b9_v_mzCDYXs[8] , 
        b9_v_mzCDYXs_4, \b9_v_mzCDYXs[9] , b9_v_mzCDYXs_3, 
        \b9_v_mzCDYXs[0] , b9_v_mzCDYXs_2, \b9_v_mzCDYXs[1] , 
        b9_v_mzCDYXs_1, \b9_v_mzCDYXs[2] , b9_v_mzCDYXs_0, 
        \b9_v_mzCDYXs[3] , b9_v_mzCDYXs, b12_2_St6KCa_jHv_8, 
        b12_2_St6KCa_jHv_7, b12_2_St6KCa_jHv_6, b12_2_St6KCa_jHv_5, 
        b12_2_St6KCa_jHv_4, b12_2_St6KCa_jHv_3, b12_2_St6KCa_jHv_2, 
        b12_2_St6KCa_jHv_1, b12_2_St6KCa_jHv_0, b12_2_St6KCa_jHv, 
        b9_v_mzCDYXs_cry_0_cy, N_24_mux, b9_v_mzCDYXs_cry_0, 
        \b9_v_mzCDYXs_RNIO1DN4_S[0] , b9_v_mzCDYXs_cry_1, 
        \b9_v_mzCDYXs_RNI4MI25_S[1] , b9_v_mzCDYXs_cry_2, 
        \b9_v_mzCDYXs_RNIHBOD5_S[2] , b9_v_mzCDYXs_cry_3, 
        \b9_v_mzCDYXs_RNIV1UO5_S[3] , b9_v_mzCDYXs_cry_4, 
        \b9_v_mzCDYXs_RNIEP346_S[4] , b9_v_mzCDYXs_cry_5, 
        \b9_v_mzCDYXs_RNIUH9F6_S[5] , b9_v_mzCDYXs_cry_6, 
        \b9_v_mzCDYXs_RNIFBFQ6_S[6] , b9_v_mzCDYXs_cry_7, 
        \b9_v_mzCDYXs_RNI16L57_S[7] , \b9_v_mzCDYXs_r_RNO_S[9] , 
        b9_v_mzCDYXs_cry_8, \b9_v_mzCDYXs_RNIK1RG7_S[8] , 
        un1_b12_2_St6KCa_jHv_s_0_462_FCO, b4_2o_z, 
        un1_b12_2_St6KCa_jHv_cry_0_net_1, un1_b12_2_St6KCa_jHv_cry_0_S, 
        un1_b12_2_St6KCa_jHv_cry_1_net_1, un1_b12_2_St6KCa_jHv_cry_1_S, 
        un1_b12_2_St6KCa_jHv_cry_2_net_1, un1_b12_2_St6KCa_jHv_cry_2_S, 
        un1_b12_2_St6KCa_jHv_cry_3_net_1, un1_b12_2_St6KCa_jHv_cry_3_S, 
        un1_b12_2_St6KCa_jHv_cry_4_net_1, un1_b12_2_St6KCa_jHv_cry_4_S, 
        un1_b12_2_St6KCa_jHv_cry_5_net_1, un1_b12_2_St6KCa_jHv_cry_5_S, 
        un1_b12_2_St6KCa_jHv_cry_6_net_1, un1_b12_2_St6KCa_jHv_cry_6_S, 
        un1_b12_2_St6KCa_jHv_cry_7_net_1, un1_b12_2_St6KCa_jHv_cry_7_S, 
        un1_b12_2_St6KCa_jHv_s_9_S, un1_b12_2_St6KCa_jHv_cry_8_net_1, 
        un1_b12_2_St6KCa_jHv_cry_8_S, b7_yYh03wy_u_0_m2_net_1, 
        un1_b13_PLF_2grFt_FH911_i_a2_0_2, \b7_nYJ_BFM_RNI3PL54[161] , 
        b8_jAA_KlCO_0_sqmuxa_4_net_1, \b7_vFW_PlM[153] , 
        \un1_b4_BVmQ[153] , \b7_vFW_PlM[113] , \un1_b4_BVmQ[113] , 
        \b7_vFW_PlM[1] , \un1_b4_BVmQ[1] , b4_ycsM, ttdo, 
        \b7_vFW_PlM[91] , \b7_vFW_PlM[61] , b3_PLF_76_net_1, 
        \b7_vFW_PlM[118] , \b7_vFW_PlM[21] , b3_PLF_74_net_1, 
        \b7_vFW_PlM[145] , \b7_vFW_PlM[83] , b3_PLF_73_net_1, 
        \b7_vFW_PlM[142] , \b7_vFW_PlM[48] , b3_PLF_72_net_1, 
        \b7_vFW_PlM[107] , \b7_vFW_PlM[77] , b3_PLF_71_net_1, 
        \b7_vFW_PlM[72] , \b7_vFW_PlM[10] , b3_PLF_70_net_1, 
        \b7_vFW_PlM[134] , \b7_vFW_PlM[37] , b3_PLF_69_net_1, 
        \b7_vFW_PlM[99] , \b7_vFW_PlM[2] , b3_PLF_68_net_1, 
        \b7_vFW_PlM[64] , \b7_vFW_PlM[15] , b3_PLF_67_net_1, 
        \b7_vFW_PlM[123] , \b7_vFW_PlM[93] , b3_PLF_66_net_1, 
        \b7_vFW_PlM[88] , \b7_vFW_PlM[26] , b3_PLF_65_net_1, 
        \b7_vFW_PlM[150] , \b7_vFW_PlM[53] , b3_PLF_64_net_1, 
        \b7_vFW_PlM[115] , \b7_vFW_PlM[18] , b3_PLF_63_net_1, 
        \b7_vFW_PlM[80] , \b7_vFW_PlM[31] , b3_PLF_62_net_1, 
        \b7_vFW_PlM[109] , \b7_vFW_PlM[12] , b3_PLF_61_net_1, 
        \b7_vFW_PlM[104] , \b7_vFW_PlM[42] , b3_PLF_60_net_1, 
        \b7_vFW_PlM[69] , \b7_vFW_PlM[7] , b3_PLF_59_net_1, 
        \b7_vFW_PlM[131] , \b7_vFW_PlM[34] , b3_PLF_58_net_1, 
        \b7_vFW_PlM[96] , \b7_vFW_PlM[47] , b3_PLF_57_net_1, 
        \b7_vFW_PlM[139] , \b7_vFW_PlM[125] , b3_PLF_56_net_1, 
        \b7_vFW_PlM[120] , \b7_vFW_PlM[58] , b3_PLF_55_net_1, 
        \b7_vFW_PlM[85] , \b7_vFW_PlM[23] , b3_PLF_54_net_1, 
        \b7_vFW_PlM[147] , \b7_vFW_PlM[50] , b3_PLF_53_net_1, 
        \b7_vFW_PlM[112] , \b7_vFW_PlM[63] , b3_PLF_52_net_1, 
        \b7_vFW_PlM[28] , \b7_vFW_PlM[14] , b3_PLF_51_net_1, 
        \b7_vFW_PlM[136] , \b7_vFW_PlM[74] , b3_PLF_50_net_1, 
        \b7_vFW_PlM[101] , \b7_vFW_PlM[39] , b3_PLF_49_net_1, 
        \b7_vFW_PlM[66] , \b7_vFW_PlM[4] , b3_PLF_48_net_1, 
        \b7_vFW_PlM[128] , \b7_vFW_PlM[79] , b3_PLF_47_net_1, 
        \b7_vFW_PlM[141] , \b7_vFW_PlM[44] , b3_PLF_46_net_1, 
        \b7_vFW_PlM[152] , \b7_vFW_PlM[90] , b3_PLF_45_net_1, 
        \b7_vFW_PlM[117] , \b7_vFW_PlM[55] , b3_PLF_44_net_1, 
        \b7_vFW_PlM[82] , \b7_vFW_PlM[20] , b3_PLF_43_net_1, 
        \b7_vFW_PlM[144] , \b7_vFW_PlM[95] , b3_PLF_42_net_1, 
        \b7_vFW_PlM[60] , \b7_vFW_PlM[30] , b3_PLF_41_net_1, 
        \b7_vFW_PlM[106] , \b7_vFW_PlM[9] , b3_PLF_40_net_1, 
        \b7_vFW_PlM[133] , \b7_vFW_PlM[71] , b3_PLF_39_net_1, 
        \b7_vFW_PlM[98] , \b7_vFW_PlM[36] , b3_PLF_38_net_1, 
        \b7_vFW_PlM[122] , \b7_vFW_PlM[76] , b3_PLF_36_net_1, 
        \b7_vFW_PlM[87] , \b7_vFW_PlM[25] , b3_PLF_35_net_1, 
        \b7_vFW_PlM[149] , \b7_vFW_PlM[52] , b3_PLF_34_net_1, 
        \b7_vFW_PlM[114] , \b7_vFW_PlM[17] , b3_PLF_33_net_1, 
        \b7_vFW_PlM[92] , \b7_vFW_PlM[62] , b3_PLF_32_net_1, 
        \b7_vFW_PlM[138] , \b7_vFW_PlM[41] , b3_PLF_31_net_1, 
        \b7_vFW_PlM[103] , \b7_vFW_PlM[6] , b3_PLF_30_net_1, 
        \b7_vFW_PlM[130] , \b7_vFW_PlM[68] , b3_PLF_29_net_1, 
        \b7_vFW_PlM[78] , \b7_vFW_PlM[33] , b3_PLF_28_net_1, 
        \b7_vFW_PlM[154] , \b7_vFW_PlM[108] , b3_PLF_27_net_1, 
        \b7_vFW_PlM[119] , \b7_vFW_PlM[57] , b3_PLF_26_net_1, 
        \b7_vFW_PlM[84] , \b7_vFW_PlM[22] , b3_PLF_25_net_1, 
        \b7_vFW_PlM[146] , \b7_vFW_PlM[49] , b3_PLF_24_net_1, 
        \b7_vFW_PlM[124] , \b7_vFW_PlM[94] , b3_PLF_23_net_1, 
        \b7_vFW_PlM[73] , \b7_vFW_PlM[11] , b3_PLF_22_net_1, 
        \b7_vFW_PlM[135] , \b7_vFW_PlM[38] , b3_PLF_21_net_1, 
        \b7_vFW_PlM[100] , \b7_vFW_PlM[3] , b3_PLF_20_net_1, 
        \b7_vFW_PlM[110] , \b7_vFW_PlM[65] , b3_PLF_19_net_1, 
        \b7_vFW_PlM[140] , \b7_vFW_PlM[27] , b3_PLF_18_net_1, 
        \b7_vFW_PlM[151] , \b7_vFW_PlM[89] , b3_PLF_17_net_1, 
        \b7_vFW_PlM[116] , \b7_vFW_PlM[54] , b3_PLF_16_net_1, 
        \b7_vFW_PlM[81] , \b7_vFW_PlM[19] , b3_PLF_15_net_1, 
        \b7_vFW_PlM[111] , \b7_vFW_PlM[13] , b3_PLF_14_net_1, 
        \b7_vFW_PlM[105] , \b7_vFW_PlM[43] , b3_PLF_13_net_1, 
        \b7_vFW_PlM[70] , \b7_vFW_PlM[8] , b3_PLF_12_net_1, 
        \b7_vFW_PlM[132] , \b7_vFW_PlM[35] , b3_PLF_11_net_1, 
        \b7_vFW_PlM[97] , \b7_vFW_PlM[0] , b3_PLF_10_net_1, 
        \b7_vFW_PlM[127] , \b7_vFW_PlM[29] , b3_PLF_9_net_1, 
        \b7_vFW_PlM[121] , \b7_vFW_PlM[59] , b3_PLF_8_net_1, 
        \b7_vFW_PlM[86] , \b7_vFW_PlM[24] , b3_PLF_7_net_1, 
        \b7_vFW_PlM[148] , \b7_vFW_PlM[51] , b3_PLF_6_net_1, 
        \b7_vFW_PlM[143] , \b7_vFW_PlM[45] , b3_PLF_4_net_1, 
        \b7_vFW_PlM[137] , \b7_vFW_PlM[75] , b3_PLF_3_net_1, 
        \b7_vFW_PlM[102] , \b7_vFW_PlM[40] , b3_PLF_2_net_1, 
        \b7_vFW_PlM[67] , \b7_vFW_PlM[5] , b3_PLF_1_net_1, 
        \b7_vFW_PlM[129] , \b7_vFW_PlM[32] , b3_PLF_0_net_1, 
        b8_jAA_KlCO_0_sqmuxa_6_net_1, m9_e_6, m9_e_5, \b7_vFW_PlM[56] , 
        b3_PLF_115_net_1, \b7_vFW_PlM[46] , b3_PLF_96_net_1, 
        \b7_vFW_PlM[16] , b3_PLF_80_net_1, \b7_vFW_PlM[126] , 
        b3_PLF_77_net_1, b8_jAA_KlCO_0_sqmuxa_8_net_1, 
        b3_PLF_134_net_1, b3_PLF_133_net_1, b3_PLF_132_net_1, 
        b3_PLF_131_net_1, b3_PLF_130_net_1, b3_PLF_129_net_1, 
        b3_PLF_128_net_1, b3_PLF_127_net_1, b3_PLF_126_net_1, 
        b3_PLF_124_net_1, b3_PLF_123_net_1, b3_PLF_122_net_1, 
        b3_PLF_121_net_1, b3_PLF_120_net_1, b3_PLF_119_net_1, 
        b3_PLF_118_net_1, b3_PLF_140_net_1, b3_PLF_136_net_1, 
        b3_PLF_135_net_1, b3_PLF_149_net_1, b3_PLF_148_net_1, 
        b3_PLF_146_net_1, b3_PLF_145_net_1, b3_PLF_151_net_1, 
        un1_b13_PLF_2grFt_FH911_i_a2_0_1, N_14_1;
    
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[6]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIFBFQ6_S[6] ), .Y(b9_v_mzCDYXs_6));
    SLE \genblk9.b7_nYJ_BFM[70]  (.D(\b7_nYJ_BFM[69] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[70] ));
    SLE \b8_FZFFLXYE[2]  (.D(\b12_2_St6KCa_jHv[2]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[2]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[102]  (.D(\b7_nYJ_BFM[101] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[102] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_6 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[6]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_5_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_6_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_6_net_1));
    SLE \genblk9.b7_nYJ_BFM[62]  (.D(\b7_nYJ_BFM[61] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[62] ));
    SLE \b12_2_St6KCa_jHv[5]  (.D(b12_2_St6KCa_jHv_4), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[5]_net_1 ));
    CFG2 #( .INIT(4'h8) )  N_406_a2_1 (.A(b10_OFWNT9khFt), .B(
        IICE_comm2iice_10), .Y(N_406_a2_1_net_1));
    SLE \genblk9.b7_nYJ_BFM[130]  (.D(\b7_nYJ_BFM[129] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[130] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_15 (.A(\b7_nYJ_BFM[82] ), .B(
        \b7_nYJ_BFM[20] ), .C(\b7_vFW_PlM[81] ), .D(\b7_vFW_PlM[19] ), 
        .Y(b3_PLF_15_net_1));
    SLE \genblk9.b7_nYJ_BFM[10]  (.D(\b7_nYJ_BFM[9] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[10] ));
    SLE \genblk9.b9_v_mzCDYXs[4]  (.D(b9_v_mzCDYXs_8), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[4] ));
    b13_vFW_xNywD_EdR_161s_10s_1024s_0s_x_0 b3_SoW (.IICE_comm2iice({
        IICE_comm2iice_11}), .b12_2_St6KCa_jHv({
        \b12_2_St6KCa_jHv[9]_net_1 , \b12_2_St6KCa_jHv[8]_net_1 , 
        \b12_2_St6KCa_jHv[7]_net_1 , \b12_2_St6KCa_jHv[6]_net_1 , 
        \b12_2_St6KCa_jHv[5]_net_1 , \b12_2_St6KCa_jHv[4]_net_1 , 
        \b12_2_St6KCa_jHv[3]_net_1 , \b12_2_St6KCa_jHv[2]_net_1 , 
        \b12_2_St6KCa_jHv[1]_net_1 , \b12_2_St6KCa_jHv[0]_net_1 }), 
        .b7_vFW_PlM({\b7_vFW_PlM[154] , \b7_vFW_PlM[153] , 
        \b7_vFW_PlM[152] , \b7_vFW_PlM[151] , \b7_vFW_PlM[150] , 
        \b7_vFW_PlM[149] , \b7_vFW_PlM[148] , \b7_vFW_PlM[147] , 
        \b7_vFW_PlM[146] , \b7_vFW_PlM[145] , \b7_vFW_PlM[144] , 
        \b7_vFW_PlM[143] , \b7_vFW_PlM[142] , \b7_vFW_PlM[141] , 
        \b7_vFW_PlM[140] , \b7_vFW_PlM[139] , \b7_vFW_PlM[138] , 
        \b7_vFW_PlM[137] , \b7_vFW_PlM[136] , \b7_vFW_PlM[135] , 
        \b7_vFW_PlM[134] , \b7_vFW_PlM[133] , \b7_vFW_PlM[132] , 
        \b7_vFW_PlM[131] , \b7_vFW_PlM[130] , \b7_vFW_PlM[129] , 
        \b7_vFW_PlM[128] , \b7_vFW_PlM[127] , \b7_vFW_PlM[126] , 
        \b7_vFW_PlM[125] , \b7_vFW_PlM[124] , \b7_vFW_PlM[123] , 
        \b7_vFW_PlM[122] , \b7_vFW_PlM[121] , \b7_vFW_PlM[120] , 
        \b7_vFW_PlM[119] , \b7_vFW_PlM[118] , \b7_vFW_PlM[117] , 
        \b7_vFW_PlM[116] , \b7_vFW_PlM[115] , \b7_vFW_PlM[114] , 
        \b7_vFW_PlM[113] , \b7_vFW_PlM[112] , \b7_vFW_PlM[111] , 
        \b7_vFW_PlM[110] , \b7_vFW_PlM[109] , \b7_vFW_PlM[108] , 
        \b7_vFW_PlM[107] , \b7_vFW_PlM[106] , \b7_vFW_PlM[105] , 
        \b7_vFW_PlM[104] , \b7_vFW_PlM[103] , \b7_vFW_PlM[102] , 
        \b7_vFW_PlM[101] , \b7_vFW_PlM[100] , \b7_vFW_PlM[99] , 
        \b7_vFW_PlM[98] , \b7_vFW_PlM[97] , \b7_vFW_PlM[96] , 
        \b7_vFW_PlM[95] , \b7_vFW_PlM[94] , \b7_vFW_PlM[93] , 
        \b7_vFW_PlM[92] , \b7_vFW_PlM[91] , \b7_vFW_PlM[90] , 
        \b7_vFW_PlM[89] , \b7_vFW_PlM[88] , \b7_vFW_PlM[87] , 
        \b7_vFW_PlM[86] , \b7_vFW_PlM[85] , \b7_vFW_PlM[84] , 
        \b7_vFW_PlM[83] , \b7_vFW_PlM[82] , \b7_vFW_PlM[81] , 
        \b7_vFW_PlM[80] , \b7_vFW_PlM[79] , \b7_vFW_PlM[78] , 
        \b7_vFW_PlM[77] , \b7_vFW_PlM[76] , \b7_vFW_PlM[75] , 
        \b7_vFW_PlM[74] , \b7_vFW_PlM[73] , \b7_vFW_PlM[72] , 
        \b7_vFW_PlM[71] , \b7_vFW_PlM[70] , \b7_vFW_PlM[69] , 
        \b7_vFW_PlM[68] , \b7_vFW_PlM[67] , \b7_vFW_PlM[66] , 
        \b7_vFW_PlM[65] , \b7_vFW_PlM[64] , \b7_vFW_PlM[63] , 
        \b7_vFW_PlM[62] , \b7_vFW_PlM[61] , \b7_vFW_PlM[60] , 
        \b7_vFW_PlM[59] , \b7_vFW_PlM[58] , \b7_vFW_PlM[57] , 
        \b7_vFW_PlM[56] , \b7_vFW_PlM[55] , \b7_vFW_PlM[54] , 
        \b7_vFW_PlM[53] , \b7_vFW_PlM[52] , \b7_vFW_PlM[51] , 
        \b7_vFW_PlM[50] , \b7_vFW_PlM[49] , \b7_vFW_PlM[48] , 
        \b7_vFW_PlM[47] , \b7_vFW_PlM[46] , \b7_vFW_PlM[45] , 
        \b7_vFW_PlM[44] , \b7_vFW_PlM[43] , \b7_vFW_PlM[42] , 
        \b7_vFW_PlM[41] , \b7_vFW_PlM[40] , \b7_vFW_PlM[39] , 
        \b7_vFW_PlM[38] , \b7_vFW_PlM[37] , \b7_vFW_PlM[36] , 
        \b7_vFW_PlM[35] , \b7_vFW_PlM[34] , \b7_vFW_PlM[33] , 
        \b7_vFW_PlM[32] , \b7_vFW_PlM[31] , \b7_vFW_PlM[30] , 
        \b7_vFW_PlM[29] , \b7_vFW_PlM[28] , \b7_vFW_PlM[27] , 
        \b7_vFW_PlM[26] , \b7_vFW_PlM[25] , \b7_vFW_PlM[24] , 
        \b7_vFW_PlM[23] , \b7_vFW_PlM[22] , \b7_vFW_PlM[21] , 
        \b7_vFW_PlM[20] , \b7_vFW_PlM[19] , \b7_vFW_PlM[18] , 
        \b7_vFW_PlM[17] , \b7_vFW_PlM[16] , \b7_vFW_PlM[15] , 
        \b7_vFW_PlM[14] , \b7_vFW_PlM[13] , \b7_vFW_PlM[12] , 
        \b7_vFW_PlM[11] , \b7_vFW_PlM[10] , \b7_vFW_PlM[9] , 
        \b7_vFW_PlM[8] , \b7_vFW_PlM[7] , \b7_vFW_PlM[6] , 
        \b7_vFW_PlM[5] , \b7_vFW_PlM[4] , \b7_vFW_PlM[3] , 
        \b7_vFW_PlM[2] , \b7_vFW_PlM[1] , \b7_vFW_PlM[0] }), 
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[154], b11_OFWNT9L_8tZ[153], 
        b11_OFWNT9L_8tZ[152], b11_OFWNT9L_8tZ[151], 
        b11_OFWNT9L_8tZ[150], b11_OFWNT9L_8tZ[149], 
        b11_OFWNT9L_8tZ[148], b11_OFWNT9L_8tZ[147], 
        b11_OFWNT9L_8tZ[146], b11_OFWNT9L_8tZ[145], 
        b11_OFWNT9L_8tZ[144], b11_OFWNT9L_8tZ[143], 
        b11_OFWNT9L_8tZ[142], b11_OFWNT9L_8tZ[141], 
        b11_OFWNT9L_8tZ[140], b11_OFWNT9L_8tZ[139], 
        b11_OFWNT9L_8tZ[138], b11_OFWNT9L_8tZ[137], 
        b11_OFWNT9L_8tZ[136], b11_OFWNT9L_8tZ[135], 
        b11_OFWNT9L_8tZ[134], b11_OFWNT9L_8tZ[133], 
        b11_OFWNT9L_8tZ[132], b11_OFWNT9L_8tZ[131], 
        b11_OFWNT9L_8tZ[130], b11_OFWNT9L_8tZ[129], 
        b11_OFWNT9L_8tZ[128], b11_OFWNT9L_8tZ[127], 
        b11_OFWNT9L_8tZ[126], b11_OFWNT9L_8tZ[125], 
        b11_OFWNT9L_8tZ[124], b11_OFWNT9L_8tZ[123], 
        b11_OFWNT9L_8tZ[122], b11_OFWNT9L_8tZ[121], 
        b11_OFWNT9L_8tZ[120], b11_OFWNT9L_8tZ[119], 
        b11_OFWNT9L_8tZ[118], b11_OFWNT9L_8tZ[117], 
        b11_OFWNT9L_8tZ[116], b11_OFWNT9L_8tZ[115], 
        b11_OFWNT9L_8tZ[114], b11_OFWNT9L_8tZ[113], 
        b11_OFWNT9L_8tZ[112], b11_OFWNT9L_8tZ[111], 
        b11_OFWNT9L_8tZ[110], b11_OFWNT9L_8tZ[109], 
        b11_OFWNT9L_8tZ[108], b11_OFWNT9L_8tZ[107], 
        b11_OFWNT9L_8tZ[106], b11_OFWNT9L_8tZ[105], 
        b11_OFWNT9L_8tZ[104], b11_OFWNT9L_8tZ[103], 
        b11_OFWNT9L_8tZ[102], b11_OFWNT9L_8tZ[101], 
        b11_OFWNT9L_8tZ[100], b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], 
        b11_OFWNT9L_8tZ[97], b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], 
        b11_OFWNT9L_8tZ[94], b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], 
        b11_OFWNT9L_8tZ[91], b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], 
        b11_OFWNT9L_8tZ[88], b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], 
        b11_OFWNT9L_8tZ[85], b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], 
        b11_OFWNT9L_8tZ[82], b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], 
        b11_OFWNT9L_8tZ[79], b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], 
        b11_OFWNT9L_8tZ[76], b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], 
        b11_OFWNT9L_8tZ[73], b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], 
        b11_OFWNT9L_8tZ[70], b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], 
        b11_OFWNT9L_8tZ[67], b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], 
        b11_OFWNT9L_8tZ[64], b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], 
        b11_OFWNT9L_8tZ[61], b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], 
        b11_OFWNT9L_8tZ[58], b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], 
        b11_OFWNT9L_8tZ[55], b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], 
        b11_OFWNT9L_8tZ[52], b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], 
        b11_OFWNT9L_8tZ[49], b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], 
        b11_OFWNT9L_8tZ[46], b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], 
        b11_OFWNT9L_8tZ[43], b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], 
        b11_OFWNT9L_8tZ[40], b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], 
        b11_OFWNT9L_8tZ[37], b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], 
        b11_OFWNT9L_8tZ[34], b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], 
        b11_OFWNT9L_8tZ[31], b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], 
        b11_OFWNT9L_8tZ[28], b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], 
        b11_OFWNT9L_8tZ[25], b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], 
        b11_OFWNT9L_8tZ[22], b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], 
        b11_OFWNT9L_8tZ[19], b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], 
        b11_OFWNT9L_8tZ[16], b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], 
        b11_OFWNT9L_8tZ[13], b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], 
        b11_OFWNT9L_8tZ[10], b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], 
        b11_OFWNT9L_8tZ[7], b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], 
        b11_OFWNT9L_8tZ[4], b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], 
        b11_OFWNT9L_8tZ[1], b11_OFWNT9L_8tZ[0]}), .b9_v_mzCDYXs_2(
        b9_v_mzCDYXs_2), .b9_v_mzCDYXs_1(b9_v_mzCDYXs_1), 
        .b9_v_mzCDYXs_0(b9_v_mzCDYXs_0), .b9_v_mzCDYXs(b9_v_mzCDYXs), 
        .b9_v_mzCDYXs_8(b9_v_mzCDYXs_8), .b9_v_mzCDYXs_7(
        b9_v_mzCDYXs_7), .b9_v_mzCDYXs_6(b9_v_mzCDYXs_6), 
        .b9_v_mzCDYXs_5(b9_v_mzCDYXs_5), .b9_v_mzCDYXs_4(
        b9_v_mzCDYXs_4), .b9_v_mzCDYXs_3(b9_v_mzCDYXs_3), .BW_clk_c(
        BW_clk_c), .b4_2o_z(b4_2o_z));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[7]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNI16L57_S[7] ), .Y(b9_v_mzCDYXs_5));
    SLE \genblk9.b7_nYJ_BFM[131]  (.D(\b7_nYJ_BFM[130] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[131] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_20 (.A(\b7_nYJ_BFM[101] ), .B(
        \b7_nYJ_BFM[4] ), .C(\b7_vFW_PlM[100] ), .D(\b7_vFW_PlM[3] ), 
        .Y(b3_PLF_20_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[8]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_8_S), .Y(b12_2_St6KCa_jHv_7));
    SLE \genblk9.b7_nYJ_BFM[40]  (.D(\b7_nYJ_BFM[39] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[40] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_3 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[3]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_2_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_3_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_3_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_55 (.A(\b7_nYJ_BFM[121] ), .B(
        \b7_nYJ_BFM[59] ), .C(\b7_vFW_PlM[120] ), .D(\b7_vFW_PlM[58] ), 
        .Y(b3_PLF_55_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[2]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_2_S), .Y(b12_2_St6KCa_jHv_1));
    SLE \genblk9.b7_nYJ_BFM[4]  (.D(\b7_nYJ_BFM[3] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[4] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[4]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIEP346_S[4] ), .Y(b9_v_mzCDYXs_8));
    SLE \genblk9.b7_nYJ_BFM[63]  (.D(\b7_nYJ_BFM[62] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[63] ));
    CFG4 #( .INIT(16'h0040) )  b12_PSyi_KyDbLbb_0_sqmuxa (.A(
        b9_PSyil9s_2_net_1), .B(b11_PSyil9s_FMZ), .C(b4_2o_z), .D(
        b8_SoWGfWYY), .Y(b12_PSyi_KyDbLbb_0_sqmuxa_net_1));
    SLE \b12_PSyi_KyDbLbb[5]  (.D(\b12_2_St6KCa_jHv[5]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[5]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[125]  (.D(\b7_nYJ_BFM[124] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[125] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_41 (.A(\b7_nYJ_BFM[61] ), .B(
        \b7_nYJ_BFM[31] ), .C(\b7_vFW_PlM[60] ), .D(\b7_vFW_PlM[30] ), 
        .Y(b3_PLF_41_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_28 (.A(\b7_nYJ_BFM[79] ), .B(
        \b7_nYJ_BFM[34] ), .C(\b7_vFW_PlM[78] ), .D(\b7_vFW_PlM[33] ), 
        .Y(b3_PLF_28_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIV1UO5[3]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[3] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_2), .S(\b9_v_mzCDYXs_RNIV1UO5_S[3] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_3));
    SLE \genblk9.b7_nYJ_BFM[80]  (.D(\b7_nYJ_BFM[79] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[80] ));
    SLE \genblk9.b7_nYJ_BFM[27]  (.D(\b7_nYJ_BFM[26] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[27] ));
    SLE \genblk9.b7_nYJ_BFM[124]  (.D(\b7_nYJ_BFM[123] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[124] ));
    SLE \genblk9.b7_nYJ_BFM[117]  (.D(\b7_nYJ_BFM[116] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[117] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_42 (.A(\b7_nYJ_BFM[145] ), .B(
        \b7_nYJ_BFM[96] ), .C(\b7_vFW_PlM[144] ), .D(\b7_vFW_PlM[95] ), 
        .Y(b3_PLF_42_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_60 (.A(\b7_nYJ_BFM[105] ), .B(
        \b7_nYJ_BFM[43] ), .C(\b7_vFW_PlM[104] ), .D(\b7_vFW_PlM[42] ), 
        .Y(b3_PLF_60_net_1));
    SLE \genblk9.b7_nYJ_BFM[72]  (.D(\b7_nYJ_BFM[71] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[72] ));
    SLE b8_jAA_KlCO (.D(VCC_net_1), .CLK(BW_clk_c), .EN(
        b8_jAA_KlCO_RNO_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        b8_jAA_KlCO_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_151 (.A(b3_PLF_123_net_1), .B(
        b3_PLF_124_net_1), .C(b3_PLF_148_net_1), .D(b3_PLF_140_net_1), 
        .Y(b3_PLF_151_net_1));
    CFG2 #( .INIT(4'hE) )  \genblk9.b7_nYJ_BFM_or[10]  (.A(
        N_406_a2_1_net_1), .B(b8_SoWGfWYY), .Y(\b7_nYJ_BFM_or[10] ));
    SLE \genblk9.b7_nYJ_BFM[66]  (.D(\b7_nYJ_BFM[65] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[66] ));
    SLE \genblk9.b7_nYJ_BFM[132]  (.D(\b7_nYJ_BFM[131] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[132] ));
    SLE \b12_PSyi_KyDbLbb[0]  (.D(\b12_2_St6KCa_jHv[0]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[0]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[4]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_4_S), .Y(b12_2_St6KCa_jHv_3));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_68 (.A(\b7_nYJ_BFM[100] ), .B(
        \b7_nYJ_BFM[3] ), .C(\b7_vFW_PlM[99] ), .D(\b7_vFW_PlM[2] ), 
        .Y(b3_PLF_68_net_1));
    SLE \genblk9.b7_nYJ_BFM[12]  (.D(\b7_nYJ_BFM[11] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[12] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNI16L57[7]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[7] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_6), .S(\b9_v_mzCDYXs_RNI16L57_S[7] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_7));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_140 (.A(b3_PLF_35_net_1), .B(
        b3_PLF_36_net_1), .C(b3_PLF_126_net_1), .D(b3_PLF_96_net_1), 
        .Y(b3_PLF_140_net_1));
    SLE \genblk9.b7_nYJ_BFM[113]  (.D(\b7_nYJ_BFM[112] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[113] ));
    SLE \genblk9.b7_nYJ_BFM[73]  (.D(\b7_nYJ_BFM[72] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[73] ));
    SLE \genblk9.b7_nYJ_BFM[61]  (.D(\b7_nYJ_BFM[60] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[61] ));
    SLE \genblk9.b7_nYJ_BFM[42]  (.D(\b7_nYJ_BFM[41] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[42] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_35 (.A(\b7_nYJ_BFM[88] ), .B(
        \b7_nYJ_BFM[26] ), .C(\b7_vFW_PlM[87] ), .D(\b7_vFW_PlM[25] ), 
        .Y(b3_PLF_35_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_2 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[2]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_1_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_2_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_2_net_1));
    SLE \b8_FZFFLXYE[6]  (.D(\b12_2_St6KCa_jHv[6]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[6]_net_1 ));
    SLE \b8_FZFFLXYE[8]  (.D(\b12_2_St6KCa_jHv[8]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[8]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_11 (.A(\b7_nYJ_BFM[133] ), .B(
        \b7_nYJ_BFM[36] ), .C(\b7_vFW_PlM[132] ), .D(\b7_vFW_PlM[35] ), 
        .Y(b3_PLF_11_net_1));
    SLE \genblk9.b7_nYJ_BFM[50]  (.D(\b7_nYJ_BFM[49] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[50] ));
    SLE \b12_PSyi_KyDbLbb[6]  (.D(\b12_2_St6KCa_jHv[6]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_71 (.A(\b7_nYJ_BFM[108] ), .B(
        \b7_nYJ_BFM[78] ), .C(\b7_vFW_PlM[107] ), .D(\b7_vFW_PlM[77] ), 
        .Y(b3_PLF_71_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[5]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIUH9F6_S[5] ), .Y(b9_v_mzCDYXs_7));
    SLE \genblk9.b7_nYJ_BFM[13]  (.D(\b7_nYJ_BFM[12] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[13] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIHBOD5[2]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[2] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_1), .S(\b9_v_mzCDYXs_RNIHBOD5_S[2] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_2));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIFBFQ6[6]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[6] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_5), .S(\b9_v_mzCDYXs_RNIFBFQ6_S[6] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_6));
    SLE \genblk9.b7_nYJ_BFM[82]  (.D(\b7_nYJ_BFM[81] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[82] ));
    SLE \genblk9.b7_nYJ_BFM[35]  (.D(\b7_nYJ_BFM[34] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[35] ));
    SLE \genblk9.b7_nYJ_BFM[119]  (.D(\b7_nYJ_BFM[118] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[119] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_12 (.A(\b7_nYJ_BFM[71] ), .B(
        \b7_nYJ_BFM[9] ), .C(\b7_vFW_PlM[70] ), .D(\b7_vFW_PlM[8] ), 
        .Y(b3_PLF_12_net_1));
    SLE \genblk9.b7_nYJ_BFM[127]  (.D(\b7_nYJ_BFM[126] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[127] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[0]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_0_S), .Y(b12_2_St6KCa_jHv));
    SLE \genblk9.b7_nYJ_BFM[24]  (.D(\b7_nYJ_BFM[23] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[24] ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_72 (.A(\b7_nYJ_BFM[143] ), .B(
        \b7_nYJ_BFM[49] ), .C(\b7_vFW_PlM[142] ), .D(\b7_vFW_PlM[48] ), 
        .Y(b3_PLF_72_net_1));
    SLE \genblk9.b7_nYJ_BFM[76]  (.D(\b7_nYJ_BFM[75] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[76] ));
    SLE \genblk9.b7_nYJ_BFM[43]  (.D(\b7_nYJ_BFM[42] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[43] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_51 (.A(\b7_nYJ_BFM[29] ), .B(
        \b7_nYJ_BFM[15] ), .C(\b7_vFW_PlM[28] ), .D(\b7_vFW_PlM[14] ), 
        .Y(b3_PLF_51_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[6]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_6_S), .Y(b12_2_St6KCa_jHv_5));
    SLE \genblk9.b7_nYJ_BFM[95]  (.D(\b7_nYJ_BFM[94] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[95] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIEP346[4]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[4] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_3), .S(\b9_v_mzCDYXs_RNIEP346_S[4] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_4));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_122 (.A(b3_PLF_26_net_1), .B(
        b3_PLF_25_net_1), .C(b3_PLF_24_net_1), .D(b3_PLF_23_net_1), .Y(
        b3_PLF_122_net_1));
    SLE \genblk9.b9_v_mzCDYXs[3]  (.D(b9_v_mzCDYXs), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[3] ));
    SLE \genblk9.b7_nYJ_BFM[29]  (.D(\b7_nYJ_BFM[28] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[29] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_52 (.A(\b7_nYJ_BFM[113] ), .B(
        \b7_nYJ_BFM[64] ), .C(\b7_vFW_PlM[112] ), .D(\b7_vFW_PlM[63] ), 
        .Y(b3_PLF_52_net_1));
    SLE \genblk9.b7_nYJ_BFM[6]  (.D(\b7_nYJ_BFM[5] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[6] ));
    SLE \genblk9.b7_nYJ_BFM[16]  (.D(\b7_nYJ_BFM[15] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[16] ));
    SLE \genblk9.b7_nYJ_BFM[83]  (.D(\b7_nYJ_BFM[82] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[83] ));
    SLE \genblk9.b7_nYJ_BFM[71]  (.D(\b7_nYJ_BFM[70] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[71] ));
    SLE \genblk9.b7_nYJ_BFM[123]  (.D(\b7_nYJ_BFM[122] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[123] ));
    SLE \genblk9.b7_nYJ_BFM[110]  (.D(\b7_nYJ_BFM[109] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[110] ));
    SLE \genblk9.b9_v_mzCDYXs[9]  (.D(b9_v_mzCDYXs_3), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[9] ));
    SLE \genblk9.b7_nYJ_BFM[46]  (.D(\b7_nYJ_BFM[45] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[46] ));
    SLE \b12_PSyi_KyDbLbb[3]  (.D(\b12_2_St6KCa_jHv[3]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_0 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[0]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_s_0_462_FCO), .S(
        un1_b12_2_St6KCa_jHv_cry_0_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIK1RG7[8]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[8] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_7), .S(\b9_v_mzCDYXs_RNIK1RG7_S[8] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_8));
    SLE \genblk9.b7_nYJ_BFM[11]  (.D(\b7_nYJ_BFM[10] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[11] ));
    SLE \genblk9.b7_nYJ_BFM[111]  (.D(\b7_nYJ_BFM[110] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[111] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_121 (.A(b3_PLF_22_net_1), .B(
        b3_PLF_21_net_1), .C(b3_PLF_20_net_1), .D(b3_PLF_19_net_1), .Y(
        b3_PLF_121_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[3]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_3_S), .Y(b12_2_St6KCa_jHv_2));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_25 (.A(\b7_nYJ_BFM[85] ), .B(
        \b7_nYJ_BFM[23] ), .C(\b7_vFW_PlM[84] ), .D(\b7_vFW_PlM[22] ), 
        .Y(b3_PLF_25_net_1));
    SLE \genblk9.b7_nYJ_BFM[52]  (.D(\b7_nYJ_BFM[51] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[52] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_s_9 (.A(VCC_net_1)
        , .B(\b12_2_St6KCa_jHv[9]_net_1 ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(un1_b12_2_St6KCa_jHv_cry_8_net_1), .S(
        un1_b12_2_St6KCa_jHv_s_9_S), .Y(), .FCO());
    SLE \genblk9.b7_nYJ_BFM[86]  (.D(\b7_nYJ_BFM[85] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[86] ));
    SLE \genblk9.b7_nYJ_BFM[41]  (.D(\b7_nYJ_BFM[40] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[41] ));
    SLE \genblk9.b7_nYJ_BFM[129]  (.D(\b7_nYJ_BFM[128] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[129] ));
    SLE \genblk9.b7_nYJ_BFM[148]  (.D(\b7_nYJ_BFM[147] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[148] ));
    SLE \genblk9.b7_nYJ_BFM[38]  (.D(\b7_nYJ_BFM[37] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[38] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_31 (.A(\b7_nYJ_BFM[139] ), .B(
        \b7_nYJ_BFM[42] ), .C(\b7_vFW_PlM[138] ), .D(\b7_vFW_PlM[41] ), 
        .Y(b3_PLF_31_net_1));
    b19_nczQ_DYg_YFaRM_oUoP_24s_1s_x_0 samplerStatus (
        .b12_PSyi_KyDbLbb({\b12_PSyi_KyDbLbb[9]_net_1 , 
        \b12_PSyi_KyDbLbb[8]_net_1 , \b12_PSyi_KyDbLbb[7]_net_1 , 
        \b12_PSyi_KyDbLbb[6]_net_1 , \b12_PSyi_KyDbLbb[5]_net_1 , 
        \b12_PSyi_KyDbLbb[4]_net_1 , \b12_PSyi_KyDbLbb[3]_net_1 , 
        \b12_PSyi_KyDbLbb[2]_net_1 , \b12_PSyi_KyDbLbb[1]_net_1 , 
        \b12_PSyi_KyDbLbb[0]_net_1 }), .b8_FZFFLXYE({
        \b8_FZFFLXYE[9]_net_1 , \b8_FZFFLXYE[8]_net_1 , 
        \b8_FZFFLXYE[7]_net_1 , \b8_FZFFLXYE[6]_net_1 , 
        \b8_FZFFLXYE[5]_net_1 , \b8_FZFFLXYE[4]_net_1 , 
        \b8_FZFFLXYE[3]_net_1 , \b8_FZFFLXYE[2]_net_1 , 
        \b8_FZFFLXYE[1]_net_1 , \b8_FZFFLXYE[0]_net_1 }), 
        .IICE_comm2iice_6(IICE_comm2iice_11), .IICE_comm2iice_4(
        IICE_comm2iice_9), .IICE_comm2iice_0(IICE_comm2iice_5), .ttdo(
        ttdo), .b8_jAA_KlCO(b8_jAA_KlCO_net_1), 
        .un1_b13_PLF_2grFt_FH911_i_a2_0_1(
        un1_b13_PLF_2grFt_FH911_i_a2_0_1), 
        .un1_b13_PLF_2grFt_FH911_i_a2_0_2(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .N_14_1(N_14_1));
    SLE \genblk9.b9_v_mzCDYXs[5]  (.D(b9_v_mzCDYXs_7), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[5] ));
    SLE \b8_FZFFLXYE[0]  (.D(\b12_2_St6KCa_jHv[0]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_s_0_462 (.A(
        VCC_net_1), .B(b4_2o_z), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(un1_b12_2_St6KCa_jHv_s_0_462_FCO));
    SLE \b12_PSyi_KyDbLbb[8]  (.D(\b12_2_St6KCa_jHv[8]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[8]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[3]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIV1UO5_S[3] ), .Y(b9_v_mzCDYXs));
    SLE \genblk9.b7_nYJ_BFM[9]  (.D(\b7_nYJ_BFM[8] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[9] ));
    SLE \genblk9.b7_nYJ_BFM[98]  (.D(\b7_nYJ_BFM[97] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[98] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_32 (.A(\b7_nYJ_BFM[93] ), .B(
        \b7_nYJ_BFM[63] ), .C(\b7_vFW_PlM[92] ), .D(\b7_vFW_PlM[62] ), 
        .Y(b3_PLF_32_net_1));
    SLE \genblk9.b7_nYJ_BFM[81]  (.D(\b7_nYJ_BFM[80] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[81] ));
    SLE \genblk9.b7_nYJ_BFM[53]  (.D(\b7_nYJ_BFM[52] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[53] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_65 (.A(\b7_nYJ_BFM[89] ), .B(
        \b7_nYJ_BFM[27] ), .C(\b7_vFW_PlM[88] ), .D(\b7_vFW_PlM[26] ), 
        .Y(b3_PLF_65_net_1));
    SLE \b8_FZFFLXYE[3]  (.D(\b12_2_St6KCa_jHv[3]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[3]_net_1 ));
    CFG4 #( .INIT(16'hFEEE) )  b3_PLF_115 (.A(\un1_b4_BVmQ[153] ), .B(
        b3_PLF_76_net_1), .C(\b7_nYJ_BFM[57] ), .D(\b7_vFW_PlM[56] ), 
        .Y(b3_PLF_115_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[1]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_1_S), .Y(b12_2_St6KCa_jHv_0));
    SLE \genblk9.b7_nYJ_BFM[112]  (.D(\b7_nYJ_BFM[111] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[112] ));
    SLE \genblk9.b7_nYJ_BFM[120]  (.D(\b7_nYJ_BFM[119] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[120] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_118 (.A(b3_PLF_10_net_1), .B(
        b3_PLF_9_net_1), .C(b3_PLF_8_net_1), .D(b3_PLF_7_net_1), .Y(
        b3_PLF_118_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_8 (.A(\b7_nYJ_BFM[122] ), .B(
        \b7_nYJ_BFM[60] ), .C(\b7_vFW_PlM[121] ), .D(\b7_vFW_PlM[59] ), 
        .Y(b3_PLF_8_net_1));
    SLE \genblk9.b7_nYJ_BFM[121]  (.D(\b7_nYJ_BFM[120] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[121] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_4 (.A(\b7_nYJ_BFM[144] ), .B(
        \b7_nYJ_BFM[46] ), .C(\b7_vFW_PlM[143] ), .D(\b7_vFW_PlM[45] ), 
        .Y(b3_PLF_4_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_128 (.A(b3_PLF_50_net_1), .B(
        b3_PLF_49_net_1), .C(b3_PLF_48_net_1), .D(b3_PLF_47_net_1), .Y(
        b3_PLF_128_net_1));
    SLE \genblk9.b7_nYJ_BFM[56]  (.D(\b7_nYJ_BFM[55] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[56] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_44 (.A(\b7_nYJ_BFM[118] ), .B(
        \b7_nYJ_BFM[56] ), .C(\b7_vFW_PlM[117] ), .D(\b7_vFW_PlM[55] ), 
        .Y(b3_PLF_44_net_1));
    SLE \genblk9.b7_nYJ_BFM[146]  (.D(\b7_nYJ_BFM[145] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[146] ));
    SLE \genblk9.b7_nYJ_BFM[65]  (.D(\b7_nYJ_BFM[64] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[65] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_46 (.A(\b7_nYJ_BFM[142] ), .B(
        \b7_nYJ_BFM[45] ), .C(\b7_vFW_PlM[141] ), .D(\b7_vFW_PlM[44] ), 
        .Y(b3_PLF_46_net_1));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b7_nYJ_BFM_RNI3PL54[161]  (.A(
        b8_nYJ_TqLY), .B(N_24_mux), .C(IICE_comm2iice_10), .D(
        b10_OFWNT9khFt), .Y(\b7_nYJ_BFM_RNI3PL54[161] ));
    CFG2 #( .INIT(4'h8) )  b8_jAA_KlCO_0_sqmuxa_4 (.A(
        \b12_2_St6KCa_jHv[7]_net_1 ), .B(\b12_2_St6KCa_jHv[8]_net_1 ), 
        .Y(b8_jAA_KlCO_0_sqmuxa_4_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_130 (.A(b3_PLF_58_net_1), .B(
        b3_PLF_57_net_1), .C(b3_PLF_56_net_1), .D(b3_PLF_55_net_1), .Y(
        b3_PLF_130_net_1));
    SLE \genblk9.b7_nYJ_BFM[51]  (.D(\b7_nYJ_BFM[50] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[51] ));
    SLE \genblk9.b7_nYJ_BFM[37]  (.D(\b7_nYJ_BFM[36] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[37] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_21 (.A(\b7_nYJ_BFM[136] ), .B(
        \b7_nYJ_BFM[39] ), .C(\b7_vFW_PlM[135] ), .D(\b7_vFW_PlM[38] ), 
        .Y(b3_PLF_21_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_126 (.A(b3_PLF_42_net_1), .B(
        b3_PLF_41_net_1), .C(b3_PLF_40_net_1), .D(b3_PLF_39_net_1), .Y(
        b3_PLF_126_net_1));
    SLE \genblk9.b7_nYJ_BFM[97]  (.D(\b7_nYJ_BFM[96] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[97] ));
    SLE \genblk9.b9_v_mzCDYXs[0]  (.D(b9_v_mzCDYXs_2), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[0] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_49 (.A(\b7_nYJ_BFM[102] ), .B(
        \b7_nYJ_BFM[40] ), .C(\b7_vFW_PlM[101] ), .D(\b7_vFW_PlM[39] ), 
        .Y(b3_PLF_49_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_5 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[5]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_4_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_5_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_5_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_22 (.A(\b7_nYJ_BFM[74] ), .B(
        \b7_nYJ_BFM[12] ), .C(\b7_vFW_PlM[73] ), .D(\b7_vFW_PlM[11] ), 
        .Y(b3_PLF_22_net_1));
    SLE \genblk9.b7_nYJ_BFM[1]  (.D(\b7_nYJ_BFM[0] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[1] ));
    SLE \genblk9.b7_nYJ_BFM[122]  (.D(\b7_nYJ_BFM[121] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[122] ));
    SLE \genblk9.b7_nYJ_BFM[20]  (.D(\b7_nYJ_BFM[19] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[20] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_47 (.A(\b7_nYJ_BFM[129] ), .B(
        \b7_nYJ_BFM[80] ), .C(\b7_vFW_PlM[128] ), .D(\b7_vFW_PlM[79] ), 
        .Y(b3_PLF_47_net_1));
    SLE \genblk9.b7_nYJ_BFM[8]  (.D(\b7_nYJ_BFM[7] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[8] ));
    SLE \genblk9.b7_nYJ_BFM[158]  (.D(\b7_nYJ_BFM[157] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[158] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_133 (.A(b3_PLF_70_net_1), .B(
        b3_PLF_69_net_1), .C(b3_PLF_68_net_1), .D(b3_PLF_67_net_1), .Y(
        b3_PLF_133_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_4 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[4]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_3_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_4_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_4_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_61 (.A(\b7_nYJ_BFM[110] ), .B(
        \b7_nYJ_BFM[13] ), .C(\b7_vFW_PlM[109] ), .D(\b7_vFW_PlM[12] ), 
        .Y(b3_PLF_61_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_1 (.A(\b7_nYJ_BFM[68] ), .B(
        \b7_nYJ_BFM[6] ), .C(\b7_vFW_PlM[67] ), .D(\b7_vFW_PlM[5] ), 
        .Y(b3_PLF_1_net_1));
    SLE \b12_PSyi_KyDbLbb[1]  (.D(\b12_2_St6KCa_jHv[1]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  b8_jAA_KlCO_0_sqmuxa (.A(
        \b12_2_St6KCa_jHv[0]_net_1 ), .B(\b12_2_St6KCa_jHv[9]_net_1 ), 
        .C(b8_jAA_KlCO_0_sqmuxa_8_net_1), .D(
        b8_jAA_KlCO_0_sqmuxa_4_net_1), .Y(b8_jAA_KlCO_0_sqmuxa_net_1));
    SLE \genblk9.b7_nYJ_BFM[75]  (.D(\b7_nYJ_BFM[74] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[75] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_14 (.A(\b7_nYJ_BFM[112] ), .B(
        \b7_nYJ_BFM[14] ), .C(\b7_vFW_PlM[111] ), .D(\b7_vFW_PlM[13] ), 
        .Y(b3_PLF_14_net_1));
    SLE \b12_PSyi_KyDbLbb[4]  (.D(\b12_2_St6KCa_jHv[4]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[4]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_134 (.A(b3_PLF_74_net_1), .B(
        b3_PLF_73_net_1), .C(b3_PLF_72_net_1), .D(b3_PLF_71_net_1), .Y(
        b3_PLF_134_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_7 (.A(\b7_nYJ_BFM[87] ), .B(
        \b7_nYJ_BFM[25] ), .C(\b7_vFW_PlM[86] ), .D(\b7_vFW_PlM[24] ), 
        .Y(b3_PLF_7_net_1));
    SLE \genblk9.b7_nYJ_BFM[108]  (.D(\b7_nYJ_BFM[107] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[108] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_16 (.A(\b7_nYJ_BFM[117] ), .B(
        \b7_nYJ_BFM[55] ), .C(\b7_vFW_PlM[116] ), .D(\b7_vFW_PlM[54] ), 
        .Y(b3_PLF_16_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_74 (.A(\b7_nYJ_BFM[119] ), .B(
        \b7_nYJ_BFM[22] ), .C(\b7_vFW_PlM[118] ), .D(\b7_vFW_PlM[21] ), 
        .Y(b3_PLF_74_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_62 (.A(\b7_nYJ_BFM[81] ), .B(
        \b7_nYJ_BFM[32] ), .C(\b7_vFW_PlM[80] ), .D(\b7_vFW_PlM[31] ), 
        .Y(b3_PLF_62_net_1));
    SLE \genblk9.b7_nYJ_BFM[160]  (.D(\b7_nYJ_BFM[159] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[160] ));
    SLE \genblk9.b7_nYJ_BFM[68]  (.D(\b7_nYJ_BFM[67] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[68] ));
    CFG4 #( .INIT(16'h2000) )  b7_yYh03wy_u_0_a2 (.A(IICE_comm2iice_0), 
        .B(IICE_comm2iice_4), .C(b7_yYh03wy_u_0_m2_net_1), .D(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .Y(b7_yYh03wy));
    SLE \b12_PSyi_KyDbLbb[2]  (.D(\b12_2_St6KCa_jHv[2]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[2]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b9_v_mzCDYXs_RNIRFPF3[7]  (.A(
        \b9_v_mzCDYXs[9] ), .B(\b9_v_mzCDYXs[7] ), .C(m9_e_6), .D(
        m9_e_5), .Y(N_24_mux));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_76 (.A(\b7_nYJ_BFM[92] ), .B(
        \b7_nYJ_BFM[62] ), .C(\b7_vFW_PlM[91] ), .D(\b7_vFW_PlM[61] ), 
        .Y(b3_PLF_76_net_1));
    SLE \genblk9.b7_nYJ_BFM[145]  (.D(\b7_nYJ_BFM[144] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[145] ));
    SLE \b12_2_St6KCa_jHv[8]  (.D(b12_2_St6KCa_jHv_7), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_1 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[1]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_0_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_1_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_1_net_1));
    SLE \genblk9.b7_nYJ_BFM[15]  (.D(\b7_nYJ_BFM[14] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[15] ));
    SLE \genblk9.b7_nYJ_BFM[144]  (.D(\b7_nYJ_BFM[143] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[144] ));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b9_v_mzCDYXs_RNIJKMC1[0]  (.A(
        \b9_v_mzCDYXs[4] ), .B(\b9_v_mzCDYXs[2] ), .C(
        \b9_v_mzCDYXs[1] ), .D(\b9_v_mzCDYXs[0] ), .Y(m9_e_6));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_54 (.A(\b7_nYJ_BFM[86] ), .B(
        \b7_nYJ_BFM[24] ), .C(\b7_vFW_PlM[85] ), .D(\b7_vFW_PlM[23] ), 
        .Y(b3_PLF_54_net_1));
    SLE \b12_PSyi_KyDbLbb[9]  (.D(\b12_2_St6KCa_jHv[9]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[9]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[161]  (.D(\b7_nYJ_BFM[160] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(b8_nYJ_TqLY));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[8]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIK1RG7_S[8] ), .Y(b9_v_mzCDYXs_4));
    SLE \genblk9.b7_nYJ_BFM[34]  (.D(\b7_nYJ_BFM[33] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[34] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_56 (.A(\b7_nYJ_BFM[140] ), .B(
        \b7_nYJ_BFM[126] ), .C(\b7_vFW_PlM[139] ), .D(
        \b7_vFW_PlM[125] ), .Y(b3_PLF_56_net_1));
    SLE \genblk9.b7_nYJ_BFM[45]  (.D(\b7_nYJ_BFM[44] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[45] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_19 (.A(\b7_nYJ_BFM[111] ), .B(
        \b7_nYJ_BFM[66] ), .C(\b7_vFW_PlM[110] ), .D(\b7_vFW_PlM[65] ), 
        .Y(b3_PLF_19_net_1));
    SLE \b12_2_St6KCa_jHv[0]  (.D(b12_2_St6KCa_jHv), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[0]_net_1 ));
    SLE \b12_PSyi_KyDbLbb[7]  (.D(\b12_2_St6KCa_jHv[7]_net_1 ), .CLK(
        BW_clk_c), .EN(b12_PSyi_KyDbLbb_0_sqmuxa_net_1), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\b12_PSyi_KyDbLbb[7]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIO1DN4[0]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[0] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_0_cy), .S(\b9_v_mzCDYXs_RNIO1DN4_S[0] )
        , .Y(), .FCO(b9_v_mzCDYXs_cry_0));
    SLE \genblk9.b7_nYJ_BFM[94]  (.D(\b7_nYJ_BFM[93] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[94] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_17 (.A(\b7_nYJ_BFM[152] ), .B(
        \b7_nYJ_BFM[90] ), .C(\b7_vFW_PlM[151] ), .D(\b7_vFW_PlM[89] ), 
        .Y(b3_PLF_17_net_1));
    SLE \b12_2_St6KCa_jHv[6]  (.D(b12_2_St6KCa_jHv_5), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[6]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[156]  (.D(\b7_nYJ_BFM[155] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[156] ));
    SLE \genblk9.b7_nYJ_BFM[39]  (.D(\b7_nYJ_BFM[38] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[39] ));
    SLE \genblk9.b7_nYJ_BFM[22]  (.D(\b7_nYJ_BFM[21] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[22] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF (.A(b3_PLF_145_net_1), .B(
        b3_PLF_151_net_1), .C(b3_PLF_149_net_1), .D(b3_PLF_146_net_1), 
        .Y(b9_OFWNT9Mxf));
    SLE \genblk9.b7_nYJ_BFM[85]  (.D(\b7_nYJ_BFM[84] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[85] ));
    CFG2 #( .INIT(4'hE) )  b8_jAA_KlCO_RNO (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .Y(
        b8_jAA_KlCO_RNO_net_1));
    CFG3 #( .INIT(8'hF8) )  b3_PLF_77 (.A(\b7_nYJ_BFM[127] ), .B(
        \b7_vFW_PlM[126] ), .C(b3_PLF_0_net_1), .Y(b3_PLF_77_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_59 (.A(\b7_nYJ_BFM[70] ), .B(
        \b7_nYJ_BFM[8] ), .C(\b7_vFW_PlM[69] ), .D(\b7_vFW_PlM[7] ), 
        .Y(b3_PLF_59_net_1));
    b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0 virOut (.IICE_comm2iice_11(
        IICE_comm2iice_11), .IICE_comm2iice_9(IICE_comm2iice_9), 
        .IICE_comm2iice_4(IICE_comm2iice_4), .IICE_comm2iice_0(
        IICE_comm2iice_0), .IICE_comm2iice_1(IICE_comm2iice_1), 
        .IICE_comm2iice_3(IICE_comm2iice_3), .IICE_comm2iice_2(
        IICE_comm2iice_2), .IICE_comm2iice_10(IICE_comm2iice_10), 
        .IICE_comm2iice_6(IICE_comm2iice_6), .IICE_comm2iice_5(
        IICE_comm2iice_5), .b4_ycsM(b4_ycsM), 
        .un1_b13_PLF_2grFt_FH911_i_a2_0_1(
        un1_b13_PLF_2grFt_FH911_i_a2_0_1), 
        .un1_b13_PLF_2grFt_FH911_i_a2_0_2(
        un1_b13_PLF_2grFt_FH911_i_a2_0_2), .N_14_1(N_14_1));
    SLE \genblk9.b9_v_mzCDYXs[8]  (.D(b9_v_mzCDYXs_4), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[8] ));
    SLE \genblk9.b7_nYJ_BFM[99]  (.D(\b7_nYJ_BFM[98] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[99] ));
    SLE \genblk9.b7_nYJ_BFM[106]  (.D(\b7_nYJ_BFM[105] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[106] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[9]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_s_9_S), .Y(b12_2_St6KCa_jHv_8));
    SLE \genblk9.b7_nYJ_BFM[78]  (.D(\b7_nYJ_BFM[77] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[78] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_57 (.A(\b7_nYJ_BFM[97] ), .B(
        \b7_nYJ_BFM[48] ), .C(\b7_vFW_PlM[96] ), .D(\b7_vFW_PlM[47] ), 
        .Y(b3_PLF_57_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_3 (.A(\b7_nYJ_BFM[138] ), .B(
        \b7_nYJ_BFM[76] ), .C(\b7_vFW_PlM[137] ), .D(\b7_vFW_PlM[75] ), 
        .Y(b3_PLF_3_net_1));
    SLE \genblk9.b7_nYJ_BFM[23]  (.D(\b7_nYJ_BFM[22] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[23] ));
    SLE \genblk9.b7_nYJ_BFM[138]  (.D(\b7_nYJ_BFM[137] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[138] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_34 (.A(\b7_nYJ_BFM[150] ), .B(
        \b7_nYJ_BFM[53] ), .C(\b7_vFW_PlM[149] ), .D(\b7_vFW_PlM[52] ), 
        .Y(b3_PLF_34_net_1));
    SLE \genblk9.b7_nYJ_BFM[67]  (.D(\b7_nYJ_BFM[66] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[67] ));
    SLE \genblk9.b7_nYJ_BFM[18]  (.D(\b7_nYJ_BFM[17] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[18] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_36 (.A(\b7_nYJ_BFM[123] ), .B(
        \b7_nYJ_BFM[77] ), .C(\b7_vFW_PlM[122] ), .D(\b7_vFW_PlM[76] ), 
        .Y(b3_PLF_36_net_1));
    SLE \genblk9.b7_nYJ_BFM[147]  (.D(\b7_nYJ_BFM[146] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[147] ));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[5]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_5_S), .Y(b12_2_St6KCa_jHv_4));
    CFG2 #( .INIT(4'h8) )  \genblk9.un1_b4_BVmQ[1]  (.A(
        \b7_vFW_PlM[1] ), .B(\b7_nYJ_BFM[2] ), .Y(\un1_b4_BVmQ[1] ));
    SLE \genblk9.b7_nYJ_BFM[48]  (.D(\b7_nYJ_BFM[47] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[48] ));
    SLE \b8_FZFFLXYE[9]  (.D(\b12_2_St6KCa_jHv[9]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[9]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_119 (.A(b3_PLF_14_net_1), .B(
        b3_PLF_13_net_1), .C(b3_PLF_12_net_1), .D(b3_PLF_11_net_1), .Y(
        b3_PLF_119_net_1));
    CFG2 #( .INIT(4'hE) )  b3_PLF_145 (.A(b3_PLF_135_net_1), .B(
        b3_PLF_136_net_1), .Y(b3_PLF_145_net_1));
    CFG2 #( .INIT(4'h8) )  \genblk9.un1_b4_BVmQ[153]  (.A(
        \b7_vFW_PlM[153] ), .B(\b7_nYJ_BFM[154] ), .Y(
        \un1_b4_BVmQ[153] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[0]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIO1DN4_S[0] ), .Y(b9_v_mzCDYXs_2));
    SLE \genblk9.b7_nYJ_BFM[55]  (.D(\b7_nYJ_BFM[54] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[55] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_43 (.A(\b7_nYJ_BFM[83] ), .B(
        \b7_nYJ_BFM[21] ), .C(\b7_vFW_PlM[82] ), .D(\b7_vFW_PlM[20] ), 
        .Y(b3_PLF_43_net_1));
    SLE b9_PSyil9s_2 (.D(b11_PSyil9s_FMZ), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(b9_PSyil9s_2_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_129 (.A(b3_PLF_54_net_1), .B(
        b3_PLF_53_net_1), .C(b3_PLF_52_net_1), .D(b3_PLF_51_net_1), .Y(
        b3_PLF_129_net_1));
    SLE \genblk9.b7_nYJ_BFM[26]  (.D(\b7_nYJ_BFM[25] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[26] ));
    SLE \b8_FZFFLXYE[4]  (.D(\b12_2_St6KCa_jHv[4]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[4]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_39 (.A(\b7_nYJ_BFM[134] ), .B(
        \b7_nYJ_BFM[72] ), .C(\b7_vFW_PlM[133] ), .D(\b7_vFW_PlM[71] ), 
        .Y(b3_PLF_39_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_148 (.A(b3_PLF_130_net_1), .B(
        b3_PLF_129_net_1), .C(b3_PLF_128_net_1), .D(b3_PLF_127_net_1), 
        .Y(b3_PLF_148_net_1));
    SLE \genblk9.b7_nYJ_BFM[88]  (.D(\b7_nYJ_BFM[87] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[88] ));
    SLE \genblk9.b7_nYJ_BFM[155]  (.D(\b7_nYJ_BFM[154] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[155] ));
    SLE \genblk9.b7_nYJ_BFM[143]  (.D(\b7_nYJ_BFM[142] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[143] ));
    SLE \genblk9.b7_nYJ_BFM[154]  (.D(\b7_nYJ_BFM[153] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[154] ));
    SLE \genblk9.b7_nYJ_BFM[21]  (.D(\b7_nYJ_BFM[20] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[21] ));
    SLE \genblk9.b7_nYJ_BFM[105]  (.D(\b7_nYJ_BFM[104] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[105] ));
    SLE \genblk9.b7_nYJ_BFM[77]  (.D(\b7_nYJ_BFM[76] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[77] ));
    SLE \genblk9.b7_nYJ_BFM[136]  (.D(\b7_nYJ_BFM[135] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[136] ));
    SLE \genblk9.b7_nYJ_BFM[104]  (.D(\b7_nYJ_BFM[103] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[104] ));
    SLE \b12_2_St6KCa_jHv[7]  (.D(b12_2_St6KCa_jHv_6), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[7]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_146 (.A(b3_PLF_122_net_1), .B(
        b3_PLF_121_net_1), .C(b3_PLF_120_net_1), .D(b3_PLF_119_net_1), 
        .Y(b3_PLF_146_net_1));
    SLE \b12_2_St6KCa_jHv[2]  (.D(b12_2_St6KCa_jHv_1), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[2]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[149]  (.D(\b7_nYJ_BFM[148] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[149] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_2 (.A(\b7_nYJ_BFM[103] ), .B(
        \b7_nYJ_BFM[41] ), .C(\b7_vFW_PlM[102] ), .D(\b7_vFW_PlM[40] ), 
        .Y(b3_PLF_2_net_1));
    SLE \genblk9.b7_nYJ_BFM[0]  (.D(b8_nYJ_TqLY), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(VCC_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[0] ));
    SLE \genblk9.b7_nYJ_BFM[64]  (.D(\b7_nYJ_BFM[63] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[64] ));
    SLE \genblk9.b7_nYJ_BFM[2]  (.D(\b7_nYJ_BFM[1] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[2] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_24 (.A(\b7_nYJ_BFM[147] ), .B(
        \b7_nYJ_BFM[50] ), .C(\b7_vFW_PlM[146] ), .D(\b7_vFW_PlM[49] ), 
        .Y(b3_PLF_24_net_1));
    ARI1 #( .INIT(20'h40040) )  \genblk9.b7_nYJ_BFM_RNIDE7C4[161]  (.A(
        b8_SoWGfWYY), .B(N_24_mux), .C(N_406_a2_1_net_1), .D(
        b8_nYJ_TqLY), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        b9_v_mzCDYXs_cry_0_cy));
    SLE \genblk9.b7_nYJ_BFM[17]  (.D(\b7_nYJ_BFM[16] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[17] ));
    SLE \b12_2_St6KCa_jHv[3]  (.D(b12_2_St6KCa_jHv_2), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_26 (.A(\b7_nYJ_BFM[120] ), .B(
        \b7_nYJ_BFM[58] ), .C(\b7_vFW_PlM[119] ), .D(\b7_vFW_PlM[57] ), 
        .Y(b3_PLF_26_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_13 (.A(\b7_nYJ_BFM[106] ), .B(
        \b7_nYJ_BFM[44] ), .C(\b7_vFW_PlM[105] ), .D(\b7_vFW_PlM[43] ), 
        .Y(b3_PLF_13_net_1));
    b11_SoWyP0zEFKY_161s_0s_6s_0s_2s_2s_0s_0s_2s_0s_x_0 b6_SoWyQD (
        .b11_OFWNT9L_8tZ({b11_OFWNT9L_8tZ[154], b11_OFWNT9L_8tZ[153], 
        b11_OFWNT9L_8tZ[152], b11_OFWNT9L_8tZ[151], 
        b11_OFWNT9L_8tZ[150], b11_OFWNT9L_8tZ[149], 
        b11_OFWNT9L_8tZ[148], b11_OFWNT9L_8tZ[147], 
        b11_OFWNT9L_8tZ[146], b11_OFWNT9L_8tZ[145], 
        b11_OFWNT9L_8tZ[144], b11_OFWNT9L_8tZ[143], 
        b11_OFWNT9L_8tZ[142], b11_OFWNT9L_8tZ[141], 
        b11_OFWNT9L_8tZ[140], b11_OFWNT9L_8tZ[139], 
        b11_OFWNT9L_8tZ[138], b11_OFWNT9L_8tZ[137], 
        b11_OFWNT9L_8tZ[136], b11_OFWNT9L_8tZ[135], 
        b11_OFWNT9L_8tZ[134], b11_OFWNT9L_8tZ[133], 
        b11_OFWNT9L_8tZ[132], b11_OFWNT9L_8tZ[131], 
        b11_OFWNT9L_8tZ[130], b11_OFWNT9L_8tZ[129], 
        b11_OFWNT9L_8tZ[128], b11_OFWNT9L_8tZ[127], 
        b11_OFWNT9L_8tZ[126], b11_OFWNT9L_8tZ[125], 
        b11_OFWNT9L_8tZ[124], b11_OFWNT9L_8tZ[123], 
        b11_OFWNT9L_8tZ[122], b11_OFWNT9L_8tZ[121], 
        b11_OFWNT9L_8tZ[120], b11_OFWNT9L_8tZ[119], 
        b11_OFWNT9L_8tZ[118], b11_OFWNT9L_8tZ[117], 
        b11_OFWNT9L_8tZ[116], b11_OFWNT9L_8tZ[115], 
        b11_OFWNT9L_8tZ[114], b11_OFWNT9L_8tZ[113], 
        b11_OFWNT9L_8tZ[112], b11_OFWNT9L_8tZ[111], 
        b11_OFWNT9L_8tZ[110], b11_OFWNT9L_8tZ[109], 
        b11_OFWNT9L_8tZ[108], b11_OFWNT9L_8tZ[107], 
        b11_OFWNT9L_8tZ[106], b11_OFWNT9L_8tZ[105], 
        b11_OFWNT9L_8tZ[104], b11_OFWNT9L_8tZ[103], 
        b11_OFWNT9L_8tZ[102], b11_OFWNT9L_8tZ[101], 
        b11_OFWNT9L_8tZ[100], b11_OFWNT9L_8tZ[99], b11_OFWNT9L_8tZ[98], 
        b11_OFWNT9L_8tZ[97], b11_OFWNT9L_8tZ[96], b11_OFWNT9L_8tZ[95], 
        b11_OFWNT9L_8tZ[94], b11_OFWNT9L_8tZ[93], b11_OFWNT9L_8tZ[92], 
        b11_OFWNT9L_8tZ[91], b11_OFWNT9L_8tZ[90], b11_OFWNT9L_8tZ[89], 
        b11_OFWNT9L_8tZ[88], b11_OFWNT9L_8tZ[87], b11_OFWNT9L_8tZ[86], 
        b11_OFWNT9L_8tZ[85], b11_OFWNT9L_8tZ[84], b11_OFWNT9L_8tZ[83], 
        b11_OFWNT9L_8tZ[82], b11_OFWNT9L_8tZ[81], b11_OFWNT9L_8tZ[80], 
        b11_OFWNT9L_8tZ[79], b11_OFWNT9L_8tZ[78], b11_OFWNT9L_8tZ[77], 
        b11_OFWNT9L_8tZ[76], b11_OFWNT9L_8tZ[75], b11_OFWNT9L_8tZ[74], 
        b11_OFWNT9L_8tZ[73], b11_OFWNT9L_8tZ[72], b11_OFWNT9L_8tZ[71], 
        b11_OFWNT9L_8tZ[70], b11_OFWNT9L_8tZ[69], b11_OFWNT9L_8tZ[68], 
        b11_OFWNT9L_8tZ[67], b11_OFWNT9L_8tZ[66], b11_OFWNT9L_8tZ[65], 
        b11_OFWNT9L_8tZ[64], b11_OFWNT9L_8tZ[63], b11_OFWNT9L_8tZ[62], 
        b11_OFWNT9L_8tZ[61], b11_OFWNT9L_8tZ[60], b11_OFWNT9L_8tZ[59], 
        b11_OFWNT9L_8tZ[58], b11_OFWNT9L_8tZ[57], b11_OFWNT9L_8tZ[56], 
        b11_OFWNT9L_8tZ[55], b11_OFWNT9L_8tZ[54], b11_OFWNT9L_8tZ[53], 
        b11_OFWNT9L_8tZ[52], b11_OFWNT9L_8tZ[51], b11_OFWNT9L_8tZ[50], 
        b11_OFWNT9L_8tZ[49], b11_OFWNT9L_8tZ[48], b11_OFWNT9L_8tZ[47], 
        b11_OFWNT9L_8tZ[46], b11_OFWNT9L_8tZ[45], b11_OFWNT9L_8tZ[44], 
        b11_OFWNT9L_8tZ[43], b11_OFWNT9L_8tZ[42], b11_OFWNT9L_8tZ[41], 
        b11_OFWNT9L_8tZ[40], b11_OFWNT9L_8tZ[39], b11_OFWNT9L_8tZ[38], 
        b11_OFWNT9L_8tZ[37], b11_OFWNT9L_8tZ[36], b11_OFWNT9L_8tZ[35], 
        b11_OFWNT9L_8tZ[34], b11_OFWNT9L_8tZ[33], b11_OFWNT9L_8tZ[32], 
        b11_OFWNT9L_8tZ[31], b11_OFWNT9L_8tZ[30], b11_OFWNT9L_8tZ[29], 
        b11_OFWNT9L_8tZ[28], b11_OFWNT9L_8tZ[27], b11_OFWNT9L_8tZ[26], 
        b11_OFWNT9L_8tZ[25], b11_OFWNT9L_8tZ[24], b11_OFWNT9L_8tZ[23], 
        b11_OFWNT9L_8tZ[22], b11_OFWNT9L_8tZ[21], b11_OFWNT9L_8tZ[20], 
        b11_OFWNT9L_8tZ[19], b11_OFWNT9L_8tZ[18], b11_OFWNT9L_8tZ[17], 
        b11_OFWNT9L_8tZ[16], b11_OFWNT9L_8tZ[15], b11_OFWNT9L_8tZ[14], 
        b11_OFWNT9L_8tZ[13], b11_OFWNT9L_8tZ[12], b11_OFWNT9L_8tZ[11], 
        b11_OFWNT9L_8tZ[10], b11_OFWNT9L_8tZ[9], b11_OFWNT9L_8tZ[8], 
        b11_OFWNT9L_8tZ[7], b11_OFWNT9L_8tZ[6], b11_OFWNT9L_8tZ[5], 
        b11_OFWNT9L_8tZ[4], b11_OFWNT9L_8tZ[3], b11_OFWNT9L_8tZ[2], 
        b11_OFWNT9L_8tZ[1], b11_OFWNT9L_8tZ[0]}), .mdiclink_reg({
        mdiclink_reg[154], mdiclink_reg[153], mdiclink_reg[152], 
        mdiclink_reg[151], mdiclink_reg[150], mdiclink_reg[149], 
        mdiclink_reg[148], mdiclink_reg[147], mdiclink_reg[146], 
        mdiclink_reg[145], mdiclink_reg[144], mdiclink_reg[143], 
        mdiclink_reg[142], mdiclink_reg[141], mdiclink_reg[140], 
        mdiclink_reg[139], mdiclink_reg[138], mdiclink_reg[137], 
        mdiclink_reg[136], mdiclink_reg[135], mdiclink_reg[134], 
        mdiclink_reg[133], mdiclink_reg[132], mdiclink_reg[131], 
        mdiclink_reg[130], mdiclink_reg[129], mdiclink_reg[128], 
        mdiclink_reg[127], mdiclink_reg[126], mdiclink_reg[125], 
        mdiclink_reg[124], mdiclink_reg[123], mdiclink_reg[122], 
        mdiclink_reg[121], mdiclink_reg[120], mdiclink_reg[119], 
        mdiclink_reg[118], mdiclink_reg[117], mdiclink_reg[116], 
        mdiclink_reg[115], mdiclink_reg[114], mdiclink_reg[113], 
        mdiclink_reg[112], mdiclink_reg[111], mdiclink_reg[110], 
        mdiclink_reg[109], mdiclink_reg[108], mdiclink_reg[107], 
        mdiclink_reg[106], mdiclink_reg[105], mdiclink_reg[104], 
        mdiclink_reg[103], mdiclink_reg[102], mdiclink_reg[101], 
        mdiclink_reg[100], mdiclink_reg[99], mdiclink_reg[98], 
        mdiclink_reg[97], mdiclink_reg[96], mdiclink_reg[95], 
        mdiclink_reg[94], mdiclink_reg[93], mdiclink_reg[92], 
        mdiclink_reg[91], mdiclink_reg[90], mdiclink_reg[89], 
        mdiclink_reg[88], mdiclink_reg[87], mdiclink_reg[86], 
        mdiclink_reg[85], mdiclink_reg[84], mdiclink_reg[83], 
        mdiclink_reg[82], mdiclink_reg[81], mdiclink_reg[80], 
        mdiclink_reg[79], mdiclink_reg[78], mdiclink_reg[77], 
        mdiclink_reg[76], mdiclink_reg[75], mdiclink_reg[74], 
        mdiclink_reg[73], mdiclink_reg[72], mdiclink_reg[71], 
        mdiclink_reg[70], mdiclink_reg[69], mdiclink_reg[68], 
        mdiclink_reg[67], mdiclink_reg[66], mdiclink_reg[65], 
        mdiclink_reg[64], mdiclink_reg[63], mdiclink_reg[62], 
        mdiclink_reg[61], mdiclink_reg[60], mdiclink_reg[59], 
        mdiclink_reg[58], mdiclink_reg[57], mdiclink_reg[56], 
        mdiclink_reg[55], mdiclink_reg[54], mdiclink_reg[53], 
        mdiclink_reg[52], mdiclink_reg[51], mdiclink_reg[50], 
        mdiclink_reg[49], mdiclink_reg[48], mdiclink_reg[47], 
        mdiclink_reg[46], mdiclink_reg[45], mdiclink_reg[44], 
        mdiclink_reg[43], mdiclink_reg[42], mdiclink_reg[41], 
        mdiclink_reg[40], mdiclink_reg[39], mdiclink_reg[38], 
        mdiclink_reg[37], mdiclink_reg[36], mdiclink_reg[35], 
        mdiclink_reg[34], mdiclink_reg[33], mdiclink_reg[32], 
        mdiclink_reg[31], mdiclink_reg[30], mdiclink_reg[29], 
        mdiclink_reg[28], mdiclink_reg[27], mdiclink_reg[26], 
        mdiclink_reg[25], mdiclink_reg[24], mdiclink_reg[23], 
        mdiclink_reg[22], mdiclink_reg[21], mdiclink_reg[20], 
        mdiclink_reg[19], mdiclink_reg[18], mdiclink_reg[17], 
        mdiclink_reg[16], mdiclink_reg[15], mdiclink_reg[14], 
        mdiclink_reg[13], mdiclink_reg[12], mdiclink_reg[11], 
        mdiclink_reg[10], mdiclink_reg[9], mdiclink_reg[8], 
        mdiclink_reg[7], mdiclink_reg[6], mdiclink_reg[5], 
        mdiclink_reg[4], mdiclink_reg[3], mdiclink_reg[2], 
        mdiclink_reg[1], mdiclink_reg[0]}), .b13_nAzGfFM_sLsv3({
        b13_nAzGfFM_sLsv3[1]}), .BW_clk_c(BW_clk_c), .b8_SoWGfWYY(
        b8_SoWGfWYY), .b4_2o_z(b4_2o_z), .b13_oRB_MqCD2_EdR_RNI9OIA(
        b13_oRB_MqCD2_EdR_RNI9OIA), .N_44(N_44));
    SLE \genblk9.b7_nYJ_BFM[47]  (.D(\b7_nYJ_BFM[46] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[47] ));
    SLE \genblk9.b9_v_mzCDYXs[7]  (.D(b9_v_mzCDYXs_5), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[7] ));
    SLE \genblk9.b7_nYJ_BFM[58]  (.D(\b7_nYJ_BFM[57] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[58] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_73 (.A(\b7_nYJ_BFM[146] ), .B(
        \b7_nYJ_BFM[84] ), .C(\b7_vFW_PlM[145] ), .D(\b7_vFW_PlM[83] ), 
        .Y(b3_PLF_73_net_1));
    SLE \genblk9.b7_nYJ_BFM[69]  (.D(\b7_nYJ_BFM[68] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[69] ));
    SLE \b8_FZFFLXYE[1]  (.D(\b12_2_St6KCa_jHv[1]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[1]_net_1 ));
    CFG4 #( .INIT(16'hFEEE) )  b3_PLF_80 (.A(\un1_b4_BVmQ[113] ), .B(
        b3_PLF_6_net_1), .C(\b7_nYJ_BFM[17] ), .D(\b7_vFW_PlM[16] ), 
        .Y(b3_PLF_80_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_132 (.A(b3_PLF_66_net_1), .B(
        b3_PLF_65_net_1), .C(b3_PLF_64_net_1), .D(b3_PLF_63_net_1), .Y(
        b3_PLF_132_net_1));
    SLE \genblk9.b7_nYJ_BFM[7]  (.D(\b7_nYJ_BFM[6] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[7] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_6 (.A(\b7_nYJ_BFM[149] ), .B(
        \b7_nYJ_BFM[52] ), .C(\b7_vFW_PlM[148] ), .D(\b7_vFW_PlM[51] ), 
        .Y(b3_PLF_6_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_40 (.A(\b7_nYJ_BFM[107] ), .B(
        \b7_nYJ_BFM[10] ), .C(\b7_vFW_PlM[106] ), .D(\b7_vFW_PlM[9] ), 
        .Y(b3_PLF_40_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_8 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[8]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_7_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_8_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_8_net_1));
    CFG2 #( .INIT(4'h8) )  \genblk9.un1_b4_BVmQ[113]  (.A(
        \b7_vFW_PlM[113] ), .B(\b7_nYJ_BFM[114] ), .Y(
        \un1_b4_BVmQ[113] ));
    SLE \genblk9.b7_nYJ_BFM[140]  (.D(\b7_nYJ_BFM[139] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[140] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_64 (.A(\b7_nYJ_BFM[151] ), .B(
        \b7_nYJ_BFM[54] ), .C(\b7_vFW_PlM[150] ), .D(\b7_vFW_PlM[53] ), 
        .Y(b3_PLF_64_net_1));
    SLE \genblk9.b7_nYJ_BFM[30]  (.D(\b7_nYJ_BFM[29] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[30] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_53 (.A(\b7_nYJ_BFM[148] ), .B(
        \b7_nYJ_BFM[51] ), .C(\b7_vFW_PlM[147] ), .D(\b7_vFW_PlM[50] ), 
        .Y(b3_PLF_53_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_29 (.A(\b7_nYJ_BFM[131] ), .B(
        \b7_nYJ_BFM[69] ), .C(\b7_vFW_PlM[130] ), .D(\b7_vFW_PlM[68] ), 
        .Y(b3_PLF_29_net_1));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[9]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_r_RNO_S[9] ), .Y(b9_v_mzCDYXs_3));
    SLE \genblk9.b7_nYJ_BFM[87]  (.D(\b7_nYJ_BFM[86] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[87] ));
    SLE \genblk9.b7_nYJ_BFM[157]  (.D(\b7_nYJ_BFM[156] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[157] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_66 (.A(\b7_nYJ_BFM[124] ), .B(
        \b7_nYJ_BFM[94] ), .C(\b7_vFW_PlM[123] ), .D(\b7_vFW_PlM[93] ), 
        .Y(b3_PLF_66_net_1));
    SLE \b8_FZFFLXYE[5]  (.D(\b12_2_St6KCa_jHv[5]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[5]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_27 (.A(\b7_nYJ_BFM[155] ), .B(
        \b7_nYJ_BFM[109] ), .C(\b7_vFW_PlM[154] ), .D(
        \b7_vFW_PlM[108] ), .Y(b3_PLF_27_net_1));
    SLE \b12_2_St6KCa_jHv[9]  (.D(b12_2_St6KCa_jHv_8), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[9]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[141]  (.D(\b7_nYJ_BFM[140] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[141] ));
    SLE \genblk9.b7_nYJ_BFM[90]  (.D(\b7_nYJ_BFM[89] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[90] ));
    CFG4 #( .INIT(16'h8000) )  b8_jAA_KlCO_0_sqmuxa_8 (.A(
        \b12_2_St6KCa_jHv[5]_net_1 ), .B(b8_jAA_KlCO_0_sqmuxa_6_net_1), 
        .C(b4_2o_z), .D(\b12_2_St6KCa_jHv[6]_net_1 ), .Y(
        b8_jAA_KlCO_0_sqmuxa_8_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_9 (.A(\b7_nYJ_BFM[128] ), .B(
        \b7_nYJ_BFM[30] ), .C(\b7_vFW_PlM[127] ), .D(\b7_vFW_PlM[29] ), 
        .Y(b3_PLF_9_net_1));
    CFG3 #( .INIT(8'h10) )  \b12_2_St6KCa_jHv_r[7]  (.A(
        b8_jAA_KlCO_0_sqmuxa_net_1), .B(b8_SoWGfWYY), .C(
        un1_b12_2_St6KCa_jHv_cry_7_S), .Y(b12_2_St6KCa_jHv_6));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_48 (.A(\b7_nYJ_BFM[67] ), .B(
        \b7_nYJ_BFM[5] ), .C(\b7_vFW_PlM[66] ), .D(\b7_vFW_PlM[4] ), 
        .Y(b3_PLF_48_net_1));
    SLE \genblk9.b7_nYJ_BFM[74]  (.D(\b7_nYJ_BFM[73] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[74] ));
    SLE \genblk9.b7_nYJ_BFM[107]  (.D(\b7_nYJ_BFM[106] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[107] ));
    SLE \genblk9.b7_nYJ_BFM[135]  (.D(\b7_nYJ_BFM[134] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[135] ));
    CFG4 #( .INIT(16'hFEEE) )  b3_PLF_96 (.A(\un1_b4_BVmQ[1] ), .B(
        b3_PLF_38_net_1), .C(\b7_nYJ_BFM[47] ), .D(\b7_vFW_PlM[46] ), 
        .Y(b3_PLF_96_net_1));
    SLE \genblk9.b7_nYJ_BFM[134]  (.D(\b7_nYJ_BFM[133] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[134] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_131 (.A(b3_PLF_62_net_1), .B(
        b3_PLF_61_net_1), .C(b3_PLF_60_net_1), .D(b3_PLF_59_net_1), .Y(
        b3_PLF_131_net_1));
    SLE \genblk9.b7_nYJ_BFM[118]  (.D(\b7_nYJ_BFM[117] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[118] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_69 (.A(\b7_nYJ_BFM[135] ), .B(
        \b7_nYJ_BFM[38] ), .C(\b7_vFW_PlM[134] ), .D(\b7_vFW_PlM[37] ), 
        .Y(b3_PLF_69_net_1));
    SLE \b8_FZFFLXYE[7]  (.D(\b12_2_St6KCa_jHv[7]_net_1 ), .CLK(
        BW_clk_c), .EN(b13_oRB_MqCD2_EdR_RNI9OIA), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b8_FZFFLXYE[7]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[153]  (.D(\b7_nYJ_BFM[152] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[153] ));
    SLE \genblk9.b7_nYJ_BFM[14]  (.D(\b7_nYJ_BFM[13] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[14] ));
    SLE \genblk9.b7_nYJ_BFM[79]  (.D(\b7_nYJ_BFM[78] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[79] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_67 (.A(\b7_nYJ_BFM[65] ), .B(
        \b7_nYJ_BFM[16] ), .C(\b7_vFW_PlM[64] ), .D(\b7_vFW_PlM[15] ), 
        .Y(b3_PLF_67_net_1));
    SLE \genblk9.b7_nYJ_BFM[44]  (.D(\b7_nYJ_BFM[43] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[44] ));
    SLE \genblk9.b7_nYJ_BFM[103]  (.D(\b7_nYJ_BFM[102] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[103] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_10 (.A(\b7_nYJ_BFM[98] ), .B(
        \b7_nYJ_BFM[1] ), .C(\b7_vFW_PlM[97] ), .D(\b7_vFW_PlM[0] ), 
        .Y(b3_PLF_10_net_1));
    SLE \genblk9.b7_nYJ_BFM[57]  (.D(\b7_nYJ_BFM[56] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[57] ));
    SLE \genblk9.b7_nYJ_BFM[19]  (.D(\b7_nYJ_BFM[18] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[19] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_33 (.A(\b7_nYJ_BFM[115] ), .B(
        \b7_nYJ_BFM[18] ), .C(\b7_vFW_PlM[114] ), .D(\b7_vFW_PlM[17] ), 
        .Y(b3_PLF_33_net_1));
    SLE \genblk9.b7_nYJ_BFM[142]  (.D(\b7_nYJ_BFM[141] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[142] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[2]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNIHBOD5_S[2] ), .Y(b9_v_mzCDYXs_0));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_70 (.A(\b7_nYJ_BFM[73] ), .B(
        \b7_nYJ_BFM[11] ), .C(\b7_vFW_PlM[72] ), .D(\b7_vFW_PlM[10] ), 
        .Y(b3_PLF_70_net_1));
    SLE \genblk9.b7_nYJ_BFM[159]  (.D(\b7_nYJ_BFM[158] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[159] ));
    SLE \genblk9.b7_nYJ_BFM[32]  (.D(\b7_nYJ_BFM[31] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[32] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_0 (.A(\b7_nYJ_BFM[130] ), .B(
        \b7_nYJ_BFM[33] ), .C(\b7_vFW_PlM[129] ), .D(\b7_vFW_PlM[32] ), 
        .Y(b3_PLF_0_net_1));
    SLE \genblk9.b7_nYJ_BFM[84]  (.D(\b7_nYJ_BFM[83] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[84] ));
    SLE \genblk9.b7_nYJ_BFM[49]  (.D(\b7_nYJ_BFM[48] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[49] ));
    SLE \genblk9.b7_nYJ_BFM[5]  (.D(\b7_nYJ_BFM[4] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[5] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_18 (.A(\b7_nYJ_BFM[141] ), .B(
        \b7_nYJ_BFM[28] ), .C(\b7_vFW_PlM[140] ), .D(\b7_vFW_PlM[27] ), 
        .Y(b3_PLF_18_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_50 (.A(\b7_nYJ_BFM[137] ), .B(
        \b7_nYJ_BFM[75] ), .C(\b7_vFW_PlM[136] ), .D(\b7_vFW_PlM[74] ), 
        .Y(b3_PLF_50_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_135 (.A(b3_PLF_2_net_1), .B(
        b3_PLF_1_net_1), .C(b3_PLF_115_net_1), .D(b3_PLF_77_net_1), .Y(
        b3_PLF_135_net_1));
    SLE \genblk9.b7_nYJ_BFM[92]  (.D(\b7_nYJ_BFM[91] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[92] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_127 (.A(b3_PLF_46_net_1), .B(
        b3_PLF_45_net_1), .C(b3_PLF_44_net_1), .D(b3_PLF_43_net_1), .Y(
        b3_PLF_127_net_1));
    SLE \b12_2_St6KCa_jHv[4]  (.D(b12_2_St6KCa_jHv_3), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNI4MI25[1]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[1] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_0), .S(\b9_v_mzCDYXs_RNI4MI25_S[1] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_1));
    SLE \genblk9.b7_nYJ_BFM[109]  (.D(\b7_nYJ_BFM[108] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[109] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_120 (.A(b3_PLF_18_net_1), .B(
        b3_PLF_17_net_1), .C(b3_PLF_16_net_1), .D(b3_PLF_15_net_1), .Y(
        b3_PLF_120_net_1));
    SLE \genblk9.b7_nYJ_BFM[116]  (.D(\b7_nYJ_BFM[115] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[116] ));
    SLE \genblk9.b7_nYJ_BFM[89]  (.D(\b7_nYJ_BFM[88] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[89] ));
    SLE \genblk9.b7_nYJ_BFM[25]  (.D(\b7_nYJ_BFM[24] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[25] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_RNIUH9F6[5]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[5] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_4), .S(\b9_v_mzCDYXs_RNIUH9F6_S[5] ), 
        .Y(), .FCO(b9_v_mzCDYXs_cry_5));
    SLE \genblk9.b7_nYJ_BFM[137]  (.D(\b7_nYJ_BFM[136] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[137] ));
    SLE \genblk9.b7_nYJ_BFM[128]  (.D(\b7_nYJ_BFM[127] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[128] ));
    SLE \genblk9.b7_nYJ_BFM[33]  (.D(\b7_nYJ_BFM[32] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[33] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_58 (.A(\b7_nYJ_BFM[132] ), .B(
        \b7_nYJ_BFM[35] ), .C(\b7_vFW_PlM[131] ), .D(\b7_vFW_PlM[34] ), 
        .Y(b3_PLF_58_net_1));
    CFG4 #( .INIT(16'h8000) )  \genblk9.b9_v_mzCDYXs_RNI24NC1[3]  (.A(
        \b9_v_mzCDYXs[8] ), .B(\b9_v_mzCDYXs[6] ), .C(
        \b9_v_mzCDYXs[5] ), .D(\b9_v_mzCDYXs[3] ), .Y(m9_e_5));
    SLE \genblk9.b7_nYJ_BFM[150]  (.D(\b7_nYJ_BFM[149] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[150] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_149 (.A(b3_PLF_134_net_1), .B(
        b3_PLF_133_net_1), .C(b3_PLF_132_net_1), .D(b3_PLF_131_net_1), 
        .Y(b3_PLF_149_net_1));
    SLE \b12_2_St6KCa_jHv[1]  (.D(b12_2_St6KCa_jHv_0), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b12_2_St6KCa_jHv[1]_net_1 ));
    SLE \genblk9.b7_nYJ_BFM[93]  (.D(\b7_nYJ_BFM[92] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[93] ));
    SLE \genblk9.b7_nYJ_BFM[3]  (.D(\b7_nYJ_BFM[2] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[3] ));
    SLE \genblk9.b7_nYJ_BFM[151]  (.D(\b7_nYJ_BFM[150] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[151] ));
    CFG3 #( .INIT(8'h10) )  \genblk9.b9_v_mzCDYXs_r[1]  (.A(
        b8_SoWGfWYY), .B(\b7_nYJ_BFM_RNI3PL54[161] ), .C(
        \b9_v_mzCDYXs_RNI4MI25_S[1] ), .Y(b9_v_mzCDYXs_1));
    SLE \genblk9.b7_nYJ_BFM[100]  (.D(\b7_nYJ_BFM[99] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[100] ));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_123 (.A(b3_PLF_30_net_1), .B(
        b3_PLF_29_net_1), .C(b3_PLF_28_net_1), .D(b3_PLF_27_net_1), .Y(
        b3_PLF_123_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_136 (.A(b3_PLF_3_net_1), .B(
        b3_PLF_4_net_1), .C(b3_PLF_118_net_1), .D(b3_PLF_80_net_1), .Y(
        b3_PLF_136_net_1));
    SLE \genblk9.b7_nYJ_BFM[60]  (.D(\b7_nYJ_BFM[59] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[60] ));
    SLE \genblk9.b9_v_mzCDYXs[1]  (.D(b9_v_mzCDYXs_1), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[1] ));
    SLE \genblk9.b7_nYJ_BFM[54]  (.D(\b7_nYJ_BFM[53] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[54] ));
    SLE \genblk9.b7_nYJ_BFM[133]  (.D(\b7_nYJ_BFM[132] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[133] ));
    SLE \genblk9.b7_nYJ_BFM[36]  (.D(\b7_nYJ_BFM[35] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[36] ));
    SLE \genblk9.b7_nYJ_BFM[101]  (.D(\b7_nYJ_BFM[100] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[101] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_23 (.A(\b7_nYJ_BFM[125] ), .B(
        \b7_nYJ_BFM[95] ), .C(\b7_vFW_PlM[124] ), .D(\b7_vFW_PlM[94] ), 
        .Y(b3_PLF_23_net_1));
    CFG3 #( .INIT(8'hE2) )  b7_yYh03wy_u_0_m2 (.A(b4_ycsM), .B(
        IICE_comm2iice_5), .C(ttdo), .Y(b7_yYh03wy_u_0_m2_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_30 (.A(\b7_nYJ_BFM[104] ), .B(
        \b7_nYJ_BFM[7] ), .C(\b7_vFW_PlM[103] ), .D(\b7_vFW_PlM[6] ), 
        .Y(b3_PLF_30_net_1));
    CFG4 #( .INIT(16'hFFFE) )  b3_PLF_124 (.A(b3_PLF_34_net_1), .B(
        b3_PLF_33_net_1), .C(b3_PLF_32_net_1), .D(b3_PLF_31_net_1), .Y(
        b3_PLF_124_net_1));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_45 (.A(\b7_nYJ_BFM[153] ), .B(
        \b7_nYJ_BFM[91] ), .C(\b7_vFW_PlM[152] ), .D(\b7_vFW_PlM[90] ), 
        .Y(b3_PLF_45_net_1));
    SLE \genblk9.b9_v_mzCDYXs[6]  (.D(b9_v_mzCDYXs_6), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[6] ));
    SLE \genblk9.b7_nYJ_BFM[96]  (.D(\b7_nYJ_BFM[95] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[96] ));
    SLE \genblk9.b7_nYJ_BFM[59]  (.D(\b7_nYJ_BFM[58] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[59] ));
    CFG4 #( .INIT(16'h8000) )  b8_jAA_KlCO_0_sqmuxa_6 (.A(
        \b12_2_St6KCa_jHv[4]_net_1 ), .B(\b12_2_St6KCa_jHv[3]_net_1 ), 
        .C(\b12_2_St6KCa_jHv[2]_net_1 ), .D(
        \b12_2_St6KCa_jHv[1]_net_1 ), .Y(b8_jAA_KlCO_0_sqmuxa_6_net_1));
    SLE \genblk9.b9_v_mzCDYXs[2]  (.D(b9_v_mzCDYXs_0), .CLK(
        IICE_comm2iice_11), .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_v_mzCDYXs[2] ));
    SLE \genblk9.b7_nYJ_BFM[31]  (.D(\b7_nYJ_BFM[30] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[31] ));
    SLE \genblk9.b7_nYJ_BFM[126]  (.D(\b7_nYJ_BFM[125] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[126] ));
    ARI1 #( .INIT(20'h4AA00) )  \genblk9.b9_v_mzCDYXs_r_RNO[9]  (.A(
        VCC_net_1), .B(\b9_v_mzCDYXs[9] ), .C(GND_net_1), .D(GND_net_1)
        , .FCI(b9_v_mzCDYXs_cry_8), .S(\b9_v_mzCDYXs_r_RNO_S[9] ), .Y()
        , .FCO());
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_38 (.A(\b7_nYJ_BFM[99] ), .B(
        \b7_nYJ_BFM[37] ), .C(\b7_vFW_PlM[98] ), .D(\b7_vFW_PlM[36] ), 
        .Y(b3_PLF_38_net_1));
    SLE \genblk9.b7_nYJ_BFM[139]  (.D(\b7_nYJ_BFM[138] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[139] ));
    SLE \genblk9.b7_nYJ_BFM[28]  (.D(\b7_nYJ_BFM[27] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[28] ));
    SLE \genblk9.b7_nYJ_BFM[152]  (.D(\b7_nYJ_BFM[151] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[152] ));
    SLE \genblk9.b7_nYJ_BFM[115]  (.D(\b7_nYJ_BFM[114] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[115] ));
    SLE \genblk9.b7_nYJ_BFM[91]  (.D(\b7_nYJ_BFM[90] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[91] ));
    CFG4 #( .INIT(16'hECA0) )  b3_PLF_63 (.A(\b7_nYJ_BFM[116] ), .B(
        \b7_nYJ_BFM[19] ), .C(\b7_vFW_PlM[115] ), .D(\b7_vFW_PlM[18] ), 
        .Y(b3_PLF_63_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_b12_2_St6KCa_jHv_cry_7 (.A(
        VCC_net_1), .B(\b12_2_St6KCa_jHv[7]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_b12_2_St6KCa_jHv_cry_6_net_1), .S(
        un1_b12_2_St6KCa_jHv_cry_7_S), .Y(), .FCO(
        un1_b12_2_St6KCa_jHv_cry_7_net_1));
    SLE \genblk9.b7_nYJ_BFM[114]  (.D(\b7_nYJ_BFM[113] ), .CLK(
        IICE_comm2iice_11), .EN(\b7_nYJ_BFM_or[10] ), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(b8_SoWGfWYY_i), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\b7_nYJ_BFM[114] ));
    
endmodule


module b7_PLF_6lN_x_0(
       b13_nvmFL_fx2rbuQ,
       N_50,
       b16_nYhI39swMeEd_A78,
       b12_vABZ3qsY_Lyh,
       b11_vABZ3qsY_XH_2,
       b15_OFWNT9khWqH_R9k,
       b12_uRrc2XfY_Lyh,
       N_48,
       b3_PLF_sn_N_17,
       b13_PSyiBgfDb_Z4D,
       b7_yYh03wy,
       b13_nUTQBgfDb_Z4D
    );
input  [6:1] b13_nvmFL_fx2rbuQ;
output N_50;
input  b16_nYhI39swMeEd_A78;
input  b12_vABZ3qsY_Lyh;
output b11_vABZ3qsY_XH_2;
input  b15_OFWNT9khWqH_R9k;
input  b12_uRrc2XfY_Lyh;
output N_48;
output b3_PLF_sn_N_17;
input  b13_PSyiBgfDb_Z4D;
input  b7_yYh03wy;
input  b13_nUTQBgfDb_Z4D;

    wire b3_PLF_sn_N_13, b3_PLF_7_bm_net_1, b3_PLF_7_am_net_1, 
        b3_PLF_sn_N_20, N_6, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hC0A0) )  b3_PLF_6 (.A(b15_OFWNT9khWqH_R9k), .B(
        b12_uRrc2XfY_Lyh), .C(b11_vABZ3qsY_XH_2), .D(
        b13_nvmFL_fx2rbuQ[3]), .Y(N_48));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h4) )  b3_PLF_sn_m14_e (.A(b13_nvmFL_fx2rbuQ[1]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .Y(b3_PLF_sn_N_20));
    CFG3 #( .INIT(8'hD8) )  b3_PLF_7_ns (.A(b3_PLF_sn_N_13), .B(
        b3_PLF_7_bm_net_1), .C(b3_PLF_7_am_net_1), .Y(N_50));
    CFG4 #( .INIT(16'h88D8) )  b3_PLF_7_bm (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(N_6), .C(b13_PSyiBgfDb_Z4D), .D(b13_nvmFL_fx2rbuQ[2]), .Y(
        b3_PLF_7_bm_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h5FFE) )  b3_PLF_sn_m16 (.A(b13_nvmFL_fx2rbuQ[6]), 
        .B(b3_PLF_sn_N_20), .C(b13_nvmFL_fx2rbuQ[5]), .D(
        b13_nvmFL_fx2rbuQ[4]), .Y(b3_PLF_sn_N_17));
    CFG3 #( .INIT(8'hD8) )  b3_PLF_7_am (.A(b13_nvmFL_fx2rbuQ[6]), .B(
        b7_yYh03wy), .C(b13_nUTQBgfDb_Z4D), .Y(b3_PLF_7_am_net_1));
    CFG3 #( .INIT(8'hE4) )  b3_PLF_0 (.A(b13_nvmFL_fx2rbuQ[1]), .B(
        b16_nYhI39swMeEd_A78), .C(b12_vABZ3qsY_Lyh), .Y(N_6));
    CFG4 #( .INIT(16'h1510) )  b3_PLF_7_ns_RNO (.A(
        b13_nvmFL_fx2rbuQ[6]), .B(b13_nvmFL_fx2rbuQ[2]), .C(
        b13_nvmFL_fx2rbuQ[3]), .D(b13_nvmFL_fx2rbuQ[1]), .Y(
        b3_PLF_sn_N_13));
    CFG3 #( .INIT(8'h01) )  b3_PLF_6_0 (.A(b13_nvmFL_fx2rbuQ[4]), .B(
        b13_nvmFL_fx2rbuQ[6]), .C(b13_nvmFL_fx2rbuQ[5]), .Y(
        b11_vABZ3qsY_XH_2));
    
endmodule


module b12_nvmFL_la1xyH_x_0(
       b13_nvmFL_fx2rbuQ,
       b11_vABZ3qsY_XH_2,
       b11_uRrc_9urXBb,
       b12_PSyiBgfDb_bd,
       b11_uRrc2XfY_XH,
       b12_PSyi2XfYF_bd,
       b12_ibScJX_E2_bd,
       b11_vABZ3qsY_XH,
       b12_nUTQBgfDb_bd,
       b15_nYhI39swMeEd_Mg,
       b14_OFWNT9khWqH_3i,
       N_48,
       b3_PLF_sn_N_17,
       N_50,
       b3_PLF
    );
input  [6:1] b13_nvmFL_fx2rbuQ;
input  b11_vABZ3qsY_XH_2;
input  b11_uRrc_9urXBb;
output b12_PSyiBgfDb_bd;
output b11_uRrc2XfY_XH;
output b12_PSyi2XfYF_bd;
output b12_ibScJX_E2_bd;
output b11_vABZ3qsY_XH;
output b12_nUTQBgfDb_bd;
output b15_nYhI39swMeEd_Mg;
output b14_OFWNT9khWqH_3i;
input  N_48;
input  b3_PLF_sn_N_17;
input  N_50;
output b3_PLF;

    wire b9_nvmFLR_ab_2, b9_nvmFLz_ab_1, b9_nvmFLp_ab_1, 
        b9_nvmFLm_ab_2_net_1, b9_nvmFLm_ab_3_net_1, GND_net_1, 
        VCC_net_1;
    
    CFG4 #( .INIT(16'h4000) )  b9_nvmFLp_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .C(b11_vABZ3qsY_XH_2), .D(
        b9_nvmFLp_ab_1), .Y(b12_PSyi2XfYF_bd));
    CFG2 #( .INIT(4'h1) )  b9_nvmFLm_ab_2 (.A(b13_nvmFL_fx2rbuQ[1]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .Y(b9_nvmFLm_ab_2_net_1));
    CFG3 #( .INIT(8'h80) )  b9_nvmFLm_ab (.A(b13_nvmFL_fx2rbuQ[4]), .B(
        b11_uRrc_9urXBb), .C(b9_nvmFLm_ab_3_net_1), .Y(
        b12_ibScJX_E2_bd));
    CFG4 #( .INIT(16'hB800) )  b3_PLF_inst_1 (.A(N_48), .B(
        b3_PLF_sn_N_17), .C(N_50), .D(b11_uRrc_9urXBb), .Y(b3_PLF));
    CFG4 #( .INIT(16'h0800) )  b9_nvmFLQ_ab (.A(b11_vABZ3qsY_XH_2), .B(
        b11_uRrc_9urXBb), .C(b13_nvmFL_fx2rbuQ[1]), .D(b9_nvmFLR_ab_2), 
        .Y(b12_nUTQBgfDb_bd));
    CFG4 #( .INIT(16'h1000) )  b9_nvmFLH_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[1]), .C(b11_vABZ3qsY_XH_2), .D(
        b9_nvmFLz_ab_1), .Y(b14_OFWNT9khWqH_3i));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h8) )  b9_nvmFLH_ab_1 (.A(b11_uRrc_9urXBb), .B(
        b13_nvmFL_fx2rbuQ[2]), .Y(b9_nvmFLz_ab_1));
    CFG2 #( .INIT(4'h8) )  b9_nvmFLR_ab_1 (.A(b11_uRrc_9urXBb), .B(
        b13_nvmFL_fx2rbuQ[1]), .Y(b9_nvmFLp_ab_1));
    CFG2 #( .INIT(4'h1) )  b9_nvmFLQ_ab_2 (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .Y(b9_nvmFLR_ab_2));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h8000) )  b9_nvmFLR_ab (.A(b11_vABZ3qsY_XH_2), .B(
        b11_uRrc_9urXBb), .C(b13_nvmFL_fx2rbuQ[1]), .D(b9_nvmFLR_ab_2), 
        .Y(b12_PSyiBgfDb_bd));
    CFG4 #( .INIT(16'h2000) )  b9_nvmFLz_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[1]), .C(b11_vABZ3qsY_XH_2), .D(
        b9_nvmFLz_ab_1), .Y(b11_uRrc2XfY_XH));
    CFG4 #( .INIT(16'h8000) )  b9_nvmFLP_ab0 (.A(b11_vABZ3qsY_XH_2), 
        .B(b11_uRrc_9urXBb), .C(b13_nvmFL_fx2rbuQ[3]), .D(
        b9_nvmFLm_ab_2_net_1), .Y(b15_nYhI39swMeEd_Mg));
    CFG4 #( .INIT(16'h2000) )  b9_nvmFLT_ab (.A(b13_nvmFL_fx2rbuQ[3]), 
        .B(b13_nvmFL_fx2rbuQ[2]), .C(b9_nvmFLp_ab_1), .D(
        b11_vABZ3qsY_XH_2), .Y(b11_vABZ3qsY_XH));
    CFG4 #( .INIT(16'h0100) )  b9_nvmFLm_ab_3 (.A(b13_nvmFL_fx2rbuQ[6])
        , .B(b13_nvmFL_fx2rbuQ[5]), .C(b13_nvmFL_fx2rbuQ[3]), .D(
        b9_nvmFLm_ab_2_net_1), .Y(b9_nvmFLm_ab_3_net_1));
    
endmodule


module b3_uKr_x(
       b13_nvmFL_fx2rbuQ,
       b11_uRrc_9urXBb,
       b3_PLy,
       b3_PLF,
       b7_PLy_PlM,
       b12_PSyiBgfDb_bd,
       b12_PSyi2XfYF_bd,
       b14_OFWNT9khWqH_3i,
       b13_PSyiBgfDb_Z4D,
       b13_PSyi2XfYF_Z4D,
       b15_OFWNT9khWqH_R9k,
       b7_yYh03wy,
       b12_nUTQBgfDb_bd,
       b11_uRrc2XfY_XH,
       b13_nUTQBgfDb_Z4D,
       b15_nYhI39swMeEd_Mg,
       b16_nYhI39swMeEd_A78,
       b11_vABZ3qsY_XH,
       b12_vABZ3qsY_Lyh,
       b12_ibScJX_E2_bd,
       b13_ibScJX_E2_Z4D,
       b12_uRrc2XfY_Lyh
    );
input  [6:1] b13_nvmFL_fx2rbuQ;
input  b11_uRrc_9urXBb;
input  b3_PLy;
output b3_PLF;
output b7_PLy_PlM;
output b12_PSyiBgfDb_bd;
output b12_PSyi2XfYF_bd;
output b14_OFWNT9khWqH_3i;
input  b13_PSyiBgfDb_Z4D;
input  b13_PSyi2XfYF_Z4D;
input  b15_OFWNT9khWqH_R9k;
input  b7_yYh03wy;
output b12_nUTQBgfDb_bd;
output b11_uRrc2XfY_XH;
input  b13_nUTQBgfDb_Z4D;
output b15_nYhI39swMeEd_Mg;
input  b16_nYhI39swMeEd_A78;
output b11_vABZ3qsY_XH;
input  b12_vABZ3qsY_Lyh;
output b12_ibScJX_E2_bd;
input  b13_ibScJX_E2_Z4D;
input  b12_uRrc2XfY_Lyh;

    wire b3_PLy_net_1, GND_net_1, VCC_net_1, \b12_PLF_6lN_8tYv.N_48 , 
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_17 , \b12_PLF_6lN_8tYv.N_50 , 
        b11_vABZ3qsY_XH_2;
    assign b3_PLy_net_1 = b3_PLy;
    assign b7_PLy_PlM = b3_PLy_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    b7_PLF_6lN_x_0 b12_PLF_6lN_8tYv (.b13_nvmFL_fx2rbuQ({
        b13_nvmFL_fx2rbuQ[6], b13_nvmFL_fx2rbuQ[5], 
        b13_nvmFL_fx2rbuQ[4], b13_nvmFL_fx2rbuQ[3], 
        b13_nvmFL_fx2rbuQ[2], b13_nvmFL_fx2rbuQ[1]}), .N_50(
        \b12_PLF_6lN_8tYv.N_50 ), .b16_nYhI39swMeEd_A78(
        b16_nYhI39swMeEd_A78), .b12_vABZ3qsY_Lyh(b12_vABZ3qsY_Lyh), 
        .b11_vABZ3qsY_XH_2(b11_vABZ3qsY_XH_2), .b15_OFWNT9khWqH_R9k(
        b15_OFWNT9khWqH_R9k), .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh), 
        .N_48(\b12_PLF_6lN_8tYv.N_48 ), .b3_PLF_sn_N_17(
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_17 ), .b13_PSyiBgfDb_Z4D(
        b13_PSyiBgfDb_Z4D), .b7_yYh03wy(b7_yYh03wy), 
        .b13_nUTQBgfDb_Z4D(b13_nUTQBgfDb_Z4D));
    b12_nvmFL_la1xyH_x_0 b10_nvscB_rGsL (.b13_nvmFL_fx2rbuQ({
        b13_nvmFL_fx2rbuQ[6], b13_nvmFL_fx2rbuQ[5], 
        b13_nvmFL_fx2rbuQ[4], b13_nvmFL_fx2rbuQ[3], 
        b13_nvmFL_fx2rbuQ[2], b13_nvmFL_fx2rbuQ[1]}), 
        .b11_vABZ3qsY_XH_2(b11_vABZ3qsY_XH_2), .b11_uRrc_9urXBb(
        b11_uRrc_9urXBb), .b12_PSyiBgfDb_bd(b12_PSyiBgfDb_bd), 
        .b11_uRrc2XfY_XH(b11_uRrc2XfY_XH), .b12_PSyi2XfYF_bd(
        b12_PSyi2XfYF_bd), .b12_ibScJX_E2_bd(b12_ibScJX_E2_bd), 
        .b11_vABZ3qsY_XH(b11_vABZ3qsY_XH), .b12_nUTQBgfDb_bd(
        b12_nUTQBgfDb_bd), .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), 
        .b14_OFWNT9khWqH_3i(b14_OFWNT9khWqH_3i), .N_48(
        \b12_PLF_6lN_8tYv.N_48 ), .b3_PLF_sn_N_17(
        \b12_PLF_6lN_8tYv.b3_PLF_sn_N_17 ), .N_50(
        \b12_PLF_6lN_8tYv.N_50 ), .b3_PLF(b3_PLF));
    
endmodule


module IICE_x(
       temp1,
       temp2,
       temp3,
       temp_count_data,
       temp_count,
       IICE_comm2iice,
       freq_1,
       freq_2,
       freq_0,
       freq_6,
       freq_10,
       freq_11,
       freq_13,
       freq_14,
       freq_15,
       BW_clk_c,
       temp_sck_c,
       temp1_csn_c,
       temp2_csn_c,
       temp3_csn_c,
       temp_so_c,
       IICE_iice2comm
    );
input  [15:0] temp1;
input  [15:0] temp2;
input  [15:0] temp3;
input  [4:0] temp_count_data;
input  [31:0] temp_count;
input  [11:0] IICE_comm2iice;
input  freq_1;
input  freq_2;
input  freq_0;
input  freq_6;
input  freq_10;
input  freq_11;
input  freq_13;
input  freq_14;
input  freq_15;
input  BW_clk_c;
input  temp_sck_c;
input  temp1_csn_c;
input  temp2_csn_c;
input  temp3_csn_c;
input  temp_so_c;
output IICE_iice2comm;

    wire \mdiclink_reg[9]_net_1 , VCC_net_1, GND_net_1, 
        \mdiclink_reg[8]_net_1 , \mdiclink_reg[7]_net_1 , 
        \mdiclink_reg[6]_net_1 , \mdiclink_reg[5]_net_1 , 
        \mdiclink_reg[4]_net_1 , \mdiclink_reg[3]_net_1 , 
        \mdiclink_reg[2]_net_1 , \mdiclink_reg[1]_net_1 , 
        \mdiclink_reg[0]_net_1 , \mdiclink_reg[24]_net_1 , 
        \mdiclink_reg[23]_net_1 , \mdiclink_reg[22]_net_1 , 
        \mdiclink_reg[21]_net_1 , \mdiclink_reg[20]_net_1 , 
        \mdiclink_reg[19]_net_1 , \mdiclink_reg[18]_net_1 , 
        \mdiclink_reg[17]_net_1 , \mdiclink_reg[16]_net_1 , 
        \mdiclink_reg[15]_net_1 , \mdiclink_reg[14]_net_1 , 
        \mdiclink_reg[13]_net_1 , \mdiclink_reg[12]_net_1 , 
        \mdiclink_reg[11]_net_1 , \mdiclink_reg[10]_net_1 , 
        \mdiclink_reg[39]_net_1 , \mdiclink_reg[38]_net_1 , 
        \mdiclink_reg[37]_net_1 , \mdiclink_reg[36]_net_1 , 
        \mdiclink_reg[35]_net_1 , \mdiclink_reg[34]_net_1 , 
        \mdiclink_reg[33]_net_1 , \mdiclink_reg[32]_net_1 , 
        \mdiclink_reg[31]_net_1 , \mdiclink_reg[30]_net_1 , 
        \mdiclink_reg[29]_net_1 , \mdiclink_reg[28]_net_1 , 
        \mdiclink_reg[27]_net_1 , \mdiclink_reg[26]_net_1 , 
        \mdiclink_reg[25]_net_1 , \mdiclink_reg[54]_net_1 , 
        \mdiclink_reg[53]_net_1 , \mdiclink_reg[52]_net_1 , 
        \mdiclink_reg[51]_net_1 , \mdiclink_reg[50]_net_1 , 
        \mdiclink_reg[49]_net_1 , \mdiclink_reg[48]_net_1 , 
        \mdiclink_reg[47]_net_1 , \mdiclink_reg[46]_net_1 , 
        \mdiclink_reg[45]_net_1 , \mdiclink_reg[44]_net_1 , 
        \mdiclink_reg[43]_net_1 , \mdiclink_reg[42]_net_1 , 
        \mdiclink_reg[41]_net_1 , \mdiclink_reg[40]_net_1 , 
        \mdiclink_reg[69]_net_1 , \mdiclink_reg[68]_net_1 , 
        \mdiclink_reg[67]_net_1 , \mdiclink_reg[66]_net_1 , 
        \mdiclink_reg[65]_net_1 , \mdiclink_reg[64]_net_1 , 
        \mdiclink_reg[63]_net_1 , \mdiclink_reg[62]_net_1 , 
        \mdiclink_reg[61]_net_1 , \mdiclink_reg[60]_net_1 , 
        \mdiclink_reg[59]_net_1 , \mdiclink_reg[58]_net_1 , 
        \mdiclink_reg[57]_net_1 , \mdiclink_reg[56]_net_1 , 
        \mdiclink_reg[55]_net_1 , \mdiclink_reg[84]_net_1 , 
        \mdiclink_reg[83]_net_1 , \mdiclink_reg[82]_net_1 , 
        \mdiclink_reg[81]_net_1 , \mdiclink_reg[80]_net_1 , 
        \mdiclink_reg[79]_net_1 , \mdiclink_reg[78]_net_1 , 
        \mdiclink_reg[77]_net_1 , \mdiclink_reg[76]_net_1 , 
        \mdiclink_reg[75]_net_1 , \mdiclink_reg[74]_net_1 , 
        \mdiclink_reg[73]_net_1 , \mdiclink_reg[72]_net_1 , 
        \mdiclink_reg[71]_net_1 , \mdiclink_reg[70]_net_1 , 
        \mdiclink_reg[99]_net_1 , \mdiclink_reg[98]_net_1 , 
        \mdiclink_reg[97]_net_1 , \mdiclink_reg[96]_net_1 , 
        \mdiclink_reg[95]_net_1 , \mdiclink_reg[94]_net_1 , 
        \mdiclink_reg[93]_net_1 , \mdiclink_reg[92]_net_1 , 
        \mdiclink_reg[91]_net_1 , \mdiclink_reg[90]_net_1 , 
        \mdiclink_reg[89]_net_1 , \mdiclink_reg[88]_net_1 , 
        \mdiclink_reg[87]_net_1 , \mdiclink_reg[86]_net_1 , 
        \mdiclink_reg[85]_net_1 , \mdiclink_reg[114]_net_1 , 
        \mdiclink_reg[113]_net_1 , \mdiclink_reg[112]_net_1 , 
        \mdiclink_reg[111]_net_1 , \mdiclink_reg[110]_net_1 , 
        \mdiclink_reg[109]_net_1 , \mdiclink_reg[108]_net_1 , 
        \mdiclink_reg[107]_net_1 , \mdiclink_reg[106]_net_1 , 
        \mdiclink_reg[105]_net_1 , \mdiclink_reg[104]_net_1 , 
        \mdiclink_reg[103]_net_1 , \mdiclink_reg[102]_net_1 , 
        \mdiclink_reg[101]_net_1 , \mdiclink_reg[100]_net_1 , 
        \mdiclink_reg[129]_net_1 , \mdiclink_reg[128]_net_1 , 
        \mdiclink_reg[127]_net_1 , \mdiclink_reg[126]_net_1 , 
        \mdiclink_reg[125]_net_1 , \mdiclink_reg[124]_net_1 , 
        \mdiclink_reg[123]_net_1 , \mdiclink_reg[122]_net_1 , 
        \mdiclink_reg[121]_net_1 , \mdiclink_reg[120]_net_1 , 
        \mdiclink_reg[119]_net_1 , \mdiclink_reg[118]_net_1 , 
        \mdiclink_reg[117]_net_1 , \mdiclink_reg[116]_net_1 , 
        \mdiclink_reg[115]_net_1 , \mdiclink_reg[144]_net_1 , 
        \mdiclink_reg[143]_net_1 , \mdiclink_reg[142]_net_1 , 
        \mdiclink_reg[141]_net_1 , \mdiclink_reg[140]_net_1 , 
        \mdiclink_reg[139]_net_1 , \mdiclink_reg[138]_net_1 , 
        \mdiclink_reg[137]_net_1 , \mdiclink_reg[136]_net_1 , 
        \mdiclink_reg[135]_net_1 , \mdiclink_reg[134]_net_1 , 
        \mdiclink_reg[133]_net_1 , \mdiclink_reg[132]_net_1 , 
        \mdiclink_reg[131]_net_1 , \mdiclink_reg[130]_net_1 , 
        \mdiclink_reg[154]_net_1 , \mdiclink_reg[153]_net_1 , 
        \mdiclink_reg[152]_net_1 , \mdiclink_reg[151]_net_1 , 
        \mdiclink_reg[150]_net_1 , \mdiclink_reg[149]_net_1 , 
        \mdiclink_reg[148]_net_1 , \mdiclink_reg[147]_net_1 , 
        \mdiclink_reg[146]_net_1 , \mdiclink_reg[145]_net_1 , b4_PLyF, 
        b8_PSyiBgYG, b8_PSyi2XYG, b10_OFWNT9khFt, b7_PSyi3wy, 
        b9_OFWNT9Mxf, b7_yYh03wy, b12_nUTQBgfDb_bd, b11_uRrc2XfY_XH, 
        b13_nUTQBgfDb_Z4D, b15_nYhI39swMeEd_Mg, b16_nYhI39swMeEd_A78, 
        b11_vABZ3qsY_XH, b12_vABZ3qsY_Lyh, b12_ibScJX_E2_bd, 
        b12_uRrc2XfY_Lyh, \b13_nAzGfFM_sLsv3[1] , \b11_OFWNT9L_8tZ[0] , 
        \b11_OFWNT9L_8tZ[1] , \b11_OFWNT9L_8tZ[2] , 
        \b11_OFWNT9L_8tZ[3] , \b11_OFWNT9L_8tZ[4] , 
        \b11_OFWNT9L_8tZ[5] , \b11_OFWNT9L_8tZ[6] , 
        \b11_OFWNT9L_8tZ[7] , \b11_OFWNT9L_8tZ[8] , 
        \b11_OFWNT9L_8tZ[9] , \b11_OFWNT9L_8tZ[10] , 
        \b11_OFWNT9L_8tZ[11] , \b11_OFWNT9L_8tZ[12] , 
        \b11_OFWNT9L_8tZ[13] , \b11_OFWNT9L_8tZ[14] , 
        \b11_OFWNT9L_8tZ[15] , \b11_OFWNT9L_8tZ[16] , 
        \b11_OFWNT9L_8tZ[17] , \b11_OFWNT9L_8tZ[18] , 
        \b11_OFWNT9L_8tZ[19] , \b11_OFWNT9L_8tZ[20] , 
        \b11_OFWNT9L_8tZ[21] , \b11_OFWNT9L_8tZ[22] , 
        \b11_OFWNT9L_8tZ[23] , \b11_OFWNT9L_8tZ[24] , 
        \b11_OFWNT9L_8tZ[25] , \b11_OFWNT9L_8tZ[26] , 
        \b11_OFWNT9L_8tZ[27] , \b11_OFWNT9L_8tZ[28] , 
        \b11_OFWNT9L_8tZ[29] , \b11_OFWNT9L_8tZ[30] , 
        \b11_OFWNT9L_8tZ[31] , \b11_OFWNT9L_8tZ[32] , 
        \b11_OFWNT9L_8tZ[33] , \b11_OFWNT9L_8tZ[34] , 
        \b11_OFWNT9L_8tZ[35] , \b11_OFWNT9L_8tZ[36] , 
        \b11_OFWNT9L_8tZ[37] , \b11_OFWNT9L_8tZ[38] , 
        \b11_OFWNT9L_8tZ[39] , \b11_OFWNT9L_8tZ[40] , 
        \b11_OFWNT9L_8tZ[41] , \b11_OFWNT9L_8tZ[42] , 
        \b11_OFWNT9L_8tZ[43] , \b11_OFWNT9L_8tZ[44] , 
        \b11_OFWNT9L_8tZ[45] , \b11_OFWNT9L_8tZ[46] , 
        \b11_OFWNT9L_8tZ[47] , \b11_OFWNT9L_8tZ[48] , 
        \b11_OFWNT9L_8tZ[49] , \b11_OFWNT9L_8tZ[50] , 
        \b11_OFWNT9L_8tZ[51] , \b11_OFWNT9L_8tZ[52] , 
        \b11_OFWNT9L_8tZ[53] , \b11_OFWNT9L_8tZ[54] , 
        \b11_OFWNT9L_8tZ[55] , \b11_OFWNT9L_8tZ[56] , 
        \b11_OFWNT9L_8tZ[57] , \b11_OFWNT9L_8tZ[58] , 
        \b11_OFWNT9L_8tZ[59] , \b11_OFWNT9L_8tZ[60] , 
        \b11_OFWNT9L_8tZ[61] , \b11_OFWNT9L_8tZ[62] , 
        \b11_OFWNT9L_8tZ[63] , \b11_OFWNT9L_8tZ[64] , 
        \b11_OFWNT9L_8tZ[65] , \b11_OFWNT9L_8tZ[66] , 
        \b11_OFWNT9L_8tZ[67] , \b11_OFWNT9L_8tZ[68] , 
        \b11_OFWNT9L_8tZ[69] , \b11_OFWNT9L_8tZ[70] , 
        \b11_OFWNT9L_8tZ[71] , \b11_OFWNT9L_8tZ[72] , 
        \b11_OFWNT9L_8tZ[73] , \b11_OFWNT9L_8tZ[74] , 
        \b11_OFWNT9L_8tZ[75] , \b11_OFWNT9L_8tZ[76] , 
        \b11_OFWNT9L_8tZ[77] , \b11_OFWNT9L_8tZ[78] , 
        \b11_OFWNT9L_8tZ[79] , \b11_OFWNT9L_8tZ[80] , 
        \b11_OFWNT9L_8tZ[81] , \b11_OFWNT9L_8tZ[82] , 
        \b11_OFWNT9L_8tZ[83] , \b11_OFWNT9L_8tZ[84] , 
        \b11_OFWNT9L_8tZ[85] , \b11_OFWNT9L_8tZ[86] , 
        \b11_OFWNT9L_8tZ[87] , \b11_OFWNT9L_8tZ[88] , 
        \b11_OFWNT9L_8tZ[89] , \b11_OFWNT9L_8tZ[90] , 
        \b11_OFWNT9L_8tZ[91] , \b11_OFWNT9L_8tZ[92] , 
        \b11_OFWNT9L_8tZ[93] , \b11_OFWNT9L_8tZ[94] , 
        \b11_OFWNT9L_8tZ[95] , \b11_OFWNT9L_8tZ[96] , 
        \b11_OFWNT9L_8tZ[97] , \b11_OFWNT9L_8tZ[98] , 
        \b11_OFWNT9L_8tZ[99] , \b11_OFWNT9L_8tZ[100] , 
        \b11_OFWNT9L_8tZ[101] , \b11_OFWNT9L_8tZ[102] , 
        \b11_OFWNT9L_8tZ[103] , \b11_OFWNT9L_8tZ[104] , 
        \b11_OFWNT9L_8tZ[105] , \b11_OFWNT9L_8tZ[106] , 
        \b11_OFWNT9L_8tZ[107] , \b11_OFWNT9L_8tZ[108] , 
        \b11_OFWNT9L_8tZ[109] , \b11_OFWNT9L_8tZ[110] , 
        \b11_OFWNT9L_8tZ[111] , \b11_OFWNT9L_8tZ[112] , 
        \b11_OFWNT9L_8tZ[113] , \b11_OFWNT9L_8tZ[114] , 
        \b11_OFWNT9L_8tZ[115] , \b11_OFWNT9L_8tZ[116] , 
        \b11_OFWNT9L_8tZ[117] , \b11_OFWNT9L_8tZ[118] , 
        \b11_OFWNT9L_8tZ[119] , \b11_OFWNT9L_8tZ[120] , 
        \b11_OFWNT9L_8tZ[121] , \b11_OFWNT9L_8tZ[122] , 
        \b11_OFWNT9L_8tZ[123] , \b11_OFWNT9L_8tZ[124] , 
        \b11_OFWNT9L_8tZ[125] , \b11_OFWNT9L_8tZ[126] , 
        \b11_OFWNT9L_8tZ[127] , \b11_OFWNT9L_8tZ[128] , 
        \b11_OFWNT9L_8tZ[129] , \b11_OFWNT9L_8tZ[130] , 
        \b11_OFWNT9L_8tZ[131] , \b11_OFWNT9L_8tZ[132] , 
        \b11_OFWNT9L_8tZ[133] , \b11_OFWNT9L_8tZ[134] , 
        \b11_OFWNT9L_8tZ[135] , \b11_OFWNT9L_8tZ[136] , 
        \b11_OFWNT9L_8tZ[137] , \b11_OFWNT9L_8tZ[138] , 
        \b11_OFWNT9L_8tZ[139] , \b11_OFWNT9L_8tZ[140] , 
        \b11_OFWNT9L_8tZ[141] , \b11_OFWNT9L_8tZ[142] , 
        \b11_OFWNT9L_8tZ[143] , \b11_OFWNT9L_8tZ[144] , 
        \b11_OFWNT9L_8tZ[145] , \b11_OFWNT9L_8tZ[146] , 
        \b11_OFWNT9L_8tZ[147] , \b11_OFWNT9L_8tZ[148] , 
        \b11_OFWNT9L_8tZ[149] , \b11_OFWNT9L_8tZ[150] , 
        \b11_OFWNT9L_8tZ[151] , \b11_OFWNT9L_8tZ[152] , 
        \b11_OFWNT9L_8tZ[153] , \b11_OFWNT9L_8tZ[154] , b8_SoWGfWYY, 
        b8_SoWGfWYY_i, N_44, b11_PSyil9s_FMZ;
    
    SLE \mdiclink_reg[89]  (.D(temp_count[26]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[89]_net_1 ));
    SLE \mdiclink_reg[117]  (.D(temp_count_data[3]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[117]_net_1 ));
    SLE \mdiclink_reg[116]  (.D(temp_count_data[4]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[116]_net_1 ));
    SLE \mdiclink_reg[110]  (.D(temp_count[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[110]_net_1 ));
    SLE \mdiclink_reg[90]  (.D(temp_count[25]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[90]_net_1 ));
    SLE \mdiclink_reg[97]  (.D(temp_count[18]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[97]_net_1 ));
    SLE \mdiclink_reg[108]  (.D(temp_count[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[108]_net_1 ));
    SLE \mdiclink_reg[134]  (.D(freq_13), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[134]_net_1 ));
    SLE \mdiclink_reg[61]  (.D(temp2[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[61]_net_1 ));
    SLE \mdiclink_reg[129]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[129]_net_1 ));
    SLE \mdiclink_reg[2]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[2]_net_1 ));
    SLE \mdiclink_reg[85]  (.D(temp_count[30]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[85]_net_1 ));
    SLE \mdiclink_reg[49]  (.D(temp1_csn_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[49]_net_1 ));
    SLE \mdiclink_reg[127]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[127]_net_1 ));
    SLE \mdiclink_reg[63]  (.D(temp2[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[63]_net_1 ));
    SLE \mdiclink_reg[126]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[126]_net_1 ));
    SLE \mdiclink_reg[120]  (.D(temp_count_data[0]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[120]_net_1 ));
    SLE \mdiclink_reg[80]  (.D(temp3[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[80]_net_1 ));
    SLE \mdiclink_reg[52]  (.D(temp2[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[52]_net_1 ));
    SLE \mdiclink_reg[87]  (.D(temp_count[28]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[87]_net_1 ));
    SLE \mdiclink_reg[68]  (.D(temp3[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[68]_net_1 ));
    SLE \mdiclink_reg[31]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[31]_net_1 ));
    SLE \mdiclink_reg[103]  (.D(temp_count[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[103]_net_1 ));
    SLE \mdiclink_reg[66]  (.D(temp2_csn_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[66]_net_1 ));
    SLE \mdiclink_reg[45]  (.D(temp1[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[45]_net_1 ));
    SLE \mdiclink_reg[54]  (.D(temp2[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[54]_net_1 ));
    SLE \mdiclink_reg[150]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[150]_net_1 ));
    SLE \mdiclink_reg[33]  (.D(temp1[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[33]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \mdiclink_reg[40]  (.D(temp1[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[40]_net_1 ));
    SLE \mdiclink_reg[105]  (.D(temp_count[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[105]_net_1 ));
    SLE \mdiclink_reg[47]  (.D(temp1[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[47]_net_1 ));
    SLE \mdiclink_reg[148]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[148]_net_1 ));
    SLE \mdiclink_reg[114]  (.D(temp_count[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[114]_net_1 ));
    SLE \mdiclink_reg[38]  (.D(temp1[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[38]_net_1 ));
    SLE \mdiclink_reg[36]  (.D(temp1[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[36]_net_1 ));
    SLE \mdiclink_reg[21]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[21]_net_1 ));
    b3_12m_x b8_12m_IFLY (.b13_nAzGfFM_sLsv3({\b13_nAzGfFM_sLsv3[1] }), 
        .IICE_comm2iice({IICE_comm2iice[11], IICE_comm2iice[10], 
        IICE_comm2iice[9], IICE_comm2iice[8]}), .mdiclink_reg({
        \mdiclink_reg[154]_net_1 , \mdiclink_reg[153]_net_1 , 
        \mdiclink_reg[152]_net_1 , \mdiclink_reg[151]_net_1 , 
        \mdiclink_reg[150]_net_1 , \mdiclink_reg[149]_net_1 , 
        \mdiclink_reg[148]_net_1 , \mdiclink_reg[147]_net_1 , 
        \mdiclink_reg[146]_net_1 , \mdiclink_reg[145]_net_1 , 
        \mdiclink_reg[144]_net_1 , \mdiclink_reg[143]_net_1 , 
        \mdiclink_reg[142]_net_1 , \mdiclink_reg[141]_net_1 , 
        \mdiclink_reg[140]_net_1 , \mdiclink_reg[139]_net_1 , 
        \mdiclink_reg[138]_net_1 , \mdiclink_reg[137]_net_1 , 
        \mdiclink_reg[136]_net_1 , \mdiclink_reg[135]_net_1 , 
        \mdiclink_reg[134]_net_1 , \mdiclink_reg[133]_net_1 , 
        \mdiclink_reg[132]_net_1 , \mdiclink_reg[131]_net_1 , 
        \mdiclink_reg[130]_net_1 , \mdiclink_reg[129]_net_1 , 
        \mdiclink_reg[128]_net_1 , \mdiclink_reg[127]_net_1 , 
        \mdiclink_reg[126]_net_1 , \mdiclink_reg[125]_net_1 , 
        \mdiclink_reg[124]_net_1 , \mdiclink_reg[123]_net_1 , 
        \mdiclink_reg[122]_net_1 , \mdiclink_reg[121]_net_1 , 
        \mdiclink_reg[120]_net_1 , \mdiclink_reg[119]_net_1 , 
        \mdiclink_reg[118]_net_1 , \mdiclink_reg[117]_net_1 , 
        \mdiclink_reg[116]_net_1 , \mdiclink_reg[115]_net_1 , 
        \mdiclink_reg[114]_net_1 , \mdiclink_reg[113]_net_1 , 
        \mdiclink_reg[112]_net_1 , \mdiclink_reg[111]_net_1 , 
        \mdiclink_reg[110]_net_1 , \mdiclink_reg[109]_net_1 , 
        \mdiclink_reg[108]_net_1 , \mdiclink_reg[107]_net_1 , 
        \mdiclink_reg[106]_net_1 , \mdiclink_reg[105]_net_1 , 
        \mdiclink_reg[104]_net_1 , \mdiclink_reg[103]_net_1 , 
        \mdiclink_reg[102]_net_1 , \mdiclink_reg[101]_net_1 , 
        \mdiclink_reg[100]_net_1 , \mdiclink_reg[99]_net_1 , 
        \mdiclink_reg[98]_net_1 , \mdiclink_reg[97]_net_1 , 
        \mdiclink_reg[96]_net_1 , \mdiclink_reg[95]_net_1 , 
        \mdiclink_reg[94]_net_1 , \mdiclink_reg[93]_net_1 , 
        \mdiclink_reg[92]_net_1 , \mdiclink_reg[91]_net_1 , 
        \mdiclink_reg[90]_net_1 , \mdiclink_reg[89]_net_1 , 
        \mdiclink_reg[88]_net_1 , \mdiclink_reg[87]_net_1 , 
        \mdiclink_reg[86]_net_1 , \mdiclink_reg[85]_net_1 , 
        \mdiclink_reg[84]_net_1 , \mdiclink_reg[83]_net_1 , 
        \mdiclink_reg[82]_net_1 , \mdiclink_reg[81]_net_1 , 
        \mdiclink_reg[80]_net_1 , \mdiclink_reg[79]_net_1 , 
        \mdiclink_reg[78]_net_1 , \mdiclink_reg[77]_net_1 , 
        \mdiclink_reg[76]_net_1 , \mdiclink_reg[75]_net_1 , 
        \mdiclink_reg[74]_net_1 , \mdiclink_reg[73]_net_1 , 
        \mdiclink_reg[72]_net_1 , \mdiclink_reg[71]_net_1 , 
        \mdiclink_reg[70]_net_1 , \mdiclink_reg[69]_net_1 , 
        \mdiclink_reg[68]_net_1 , \mdiclink_reg[67]_net_1 , 
        \mdiclink_reg[66]_net_1 , \mdiclink_reg[65]_net_1 , 
        \mdiclink_reg[64]_net_1 , \mdiclink_reg[63]_net_1 , 
        \mdiclink_reg[62]_net_1 , \mdiclink_reg[61]_net_1 , 
        \mdiclink_reg[60]_net_1 , \mdiclink_reg[59]_net_1 , 
        \mdiclink_reg[58]_net_1 , \mdiclink_reg[57]_net_1 , 
        \mdiclink_reg[56]_net_1 , \mdiclink_reg[55]_net_1 , 
        \mdiclink_reg[54]_net_1 , \mdiclink_reg[53]_net_1 , 
        \mdiclink_reg[52]_net_1 , \mdiclink_reg[51]_net_1 , 
        \mdiclink_reg[50]_net_1 , \mdiclink_reg[49]_net_1 , 
        \mdiclink_reg[48]_net_1 , \mdiclink_reg[47]_net_1 , 
        \mdiclink_reg[46]_net_1 , \mdiclink_reg[45]_net_1 , 
        \mdiclink_reg[44]_net_1 , \mdiclink_reg[43]_net_1 , 
        \mdiclink_reg[42]_net_1 , \mdiclink_reg[41]_net_1 , 
        \mdiclink_reg[40]_net_1 , \mdiclink_reg[39]_net_1 , 
        \mdiclink_reg[38]_net_1 , \mdiclink_reg[37]_net_1 , 
        \mdiclink_reg[36]_net_1 , \mdiclink_reg[35]_net_1 , 
        \mdiclink_reg[34]_net_1 , \mdiclink_reg[33]_net_1 , 
        \mdiclink_reg[32]_net_1 , \mdiclink_reg[31]_net_1 , 
        \mdiclink_reg[30]_net_1 , \mdiclink_reg[29]_net_1 , 
        \mdiclink_reg[28]_net_1 , \mdiclink_reg[27]_net_1 , 
        \mdiclink_reg[26]_net_1 , \mdiclink_reg[25]_net_1 , 
        \mdiclink_reg[24]_net_1 , \mdiclink_reg[23]_net_1 , 
        \mdiclink_reg[22]_net_1 , \mdiclink_reg[21]_net_1 , 
        \mdiclink_reg[20]_net_1 , \mdiclink_reg[19]_net_1 , 
        \mdiclink_reg[18]_net_1 , \mdiclink_reg[17]_net_1 , 
        \mdiclink_reg[16]_net_1 , \mdiclink_reg[15]_net_1 , 
        \mdiclink_reg[14]_net_1 , \mdiclink_reg[13]_net_1 , 
        \mdiclink_reg[12]_net_1 , \mdiclink_reg[11]_net_1 , 
        \mdiclink_reg[10]_net_1 , \mdiclink_reg[9]_net_1 , 
        \mdiclink_reg[8]_net_1 , \mdiclink_reg[7]_net_1 , 
        \mdiclink_reg[6]_net_1 , \mdiclink_reg[5]_net_1 , 
        \mdiclink_reg[4]_net_1 , \mdiclink_reg[3]_net_1 , 
        \mdiclink_reg[2]_net_1 , \mdiclink_reg[1]_net_1 , 
        \mdiclink_reg[0]_net_1 }), .b11_OFWNT9L_8tZ({
        \b11_OFWNT9L_8tZ[154] , \b11_OFWNT9L_8tZ[153] , 
        \b11_OFWNT9L_8tZ[152] , \b11_OFWNT9L_8tZ[151] , 
        \b11_OFWNT9L_8tZ[150] , \b11_OFWNT9L_8tZ[149] , 
        \b11_OFWNT9L_8tZ[148] , \b11_OFWNT9L_8tZ[147] , 
        \b11_OFWNT9L_8tZ[146] , \b11_OFWNT9L_8tZ[145] , 
        \b11_OFWNT9L_8tZ[144] , \b11_OFWNT9L_8tZ[143] , 
        \b11_OFWNT9L_8tZ[142] , \b11_OFWNT9L_8tZ[141] , 
        \b11_OFWNT9L_8tZ[140] , \b11_OFWNT9L_8tZ[139] , 
        \b11_OFWNT9L_8tZ[138] , \b11_OFWNT9L_8tZ[137] , 
        \b11_OFWNT9L_8tZ[136] , \b11_OFWNT9L_8tZ[135] , 
        \b11_OFWNT9L_8tZ[134] , \b11_OFWNT9L_8tZ[133] , 
        \b11_OFWNT9L_8tZ[132] , \b11_OFWNT9L_8tZ[131] , 
        \b11_OFWNT9L_8tZ[130] , \b11_OFWNT9L_8tZ[129] , 
        \b11_OFWNT9L_8tZ[128] , \b11_OFWNT9L_8tZ[127] , 
        \b11_OFWNT9L_8tZ[126] , \b11_OFWNT9L_8tZ[125] , 
        \b11_OFWNT9L_8tZ[124] , \b11_OFWNT9L_8tZ[123] , 
        \b11_OFWNT9L_8tZ[122] , \b11_OFWNT9L_8tZ[121] , 
        \b11_OFWNT9L_8tZ[120] , \b11_OFWNT9L_8tZ[119] , 
        \b11_OFWNT9L_8tZ[118] , \b11_OFWNT9L_8tZ[117] , 
        \b11_OFWNT9L_8tZ[116] , \b11_OFWNT9L_8tZ[115] , 
        \b11_OFWNT9L_8tZ[114] , \b11_OFWNT9L_8tZ[113] , 
        \b11_OFWNT9L_8tZ[112] , \b11_OFWNT9L_8tZ[111] , 
        \b11_OFWNT9L_8tZ[110] , \b11_OFWNT9L_8tZ[109] , 
        \b11_OFWNT9L_8tZ[108] , \b11_OFWNT9L_8tZ[107] , 
        \b11_OFWNT9L_8tZ[106] , \b11_OFWNT9L_8tZ[105] , 
        \b11_OFWNT9L_8tZ[104] , \b11_OFWNT9L_8tZ[103] , 
        \b11_OFWNT9L_8tZ[102] , \b11_OFWNT9L_8tZ[101] , 
        \b11_OFWNT9L_8tZ[100] , \b11_OFWNT9L_8tZ[99] , 
        \b11_OFWNT9L_8tZ[98] , \b11_OFWNT9L_8tZ[97] , 
        \b11_OFWNT9L_8tZ[96] , \b11_OFWNT9L_8tZ[95] , 
        \b11_OFWNT9L_8tZ[94] , \b11_OFWNT9L_8tZ[93] , 
        \b11_OFWNT9L_8tZ[92] , \b11_OFWNT9L_8tZ[91] , 
        \b11_OFWNT9L_8tZ[90] , \b11_OFWNT9L_8tZ[89] , 
        \b11_OFWNT9L_8tZ[88] , \b11_OFWNT9L_8tZ[87] , 
        \b11_OFWNT9L_8tZ[86] , \b11_OFWNT9L_8tZ[85] , 
        \b11_OFWNT9L_8tZ[84] , \b11_OFWNT9L_8tZ[83] , 
        \b11_OFWNT9L_8tZ[82] , \b11_OFWNT9L_8tZ[81] , 
        \b11_OFWNT9L_8tZ[80] , \b11_OFWNT9L_8tZ[79] , 
        \b11_OFWNT9L_8tZ[78] , \b11_OFWNT9L_8tZ[77] , 
        \b11_OFWNT9L_8tZ[76] , \b11_OFWNT9L_8tZ[75] , 
        \b11_OFWNT9L_8tZ[74] , \b11_OFWNT9L_8tZ[73] , 
        \b11_OFWNT9L_8tZ[72] , \b11_OFWNT9L_8tZ[71] , 
        \b11_OFWNT9L_8tZ[70] , \b11_OFWNT9L_8tZ[69] , 
        \b11_OFWNT9L_8tZ[68] , \b11_OFWNT9L_8tZ[67] , 
        \b11_OFWNT9L_8tZ[66] , \b11_OFWNT9L_8tZ[65] , 
        \b11_OFWNT9L_8tZ[64] , \b11_OFWNT9L_8tZ[63] , 
        \b11_OFWNT9L_8tZ[62] , \b11_OFWNT9L_8tZ[61] , 
        \b11_OFWNT9L_8tZ[60] , \b11_OFWNT9L_8tZ[59] , 
        \b11_OFWNT9L_8tZ[58] , \b11_OFWNT9L_8tZ[57] , 
        \b11_OFWNT9L_8tZ[56] , \b11_OFWNT9L_8tZ[55] , 
        \b11_OFWNT9L_8tZ[54] , \b11_OFWNT9L_8tZ[53] , 
        \b11_OFWNT9L_8tZ[52] , \b11_OFWNT9L_8tZ[51] , 
        \b11_OFWNT9L_8tZ[50] , \b11_OFWNT9L_8tZ[49] , 
        \b11_OFWNT9L_8tZ[48] , \b11_OFWNT9L_8tZ[47] , 
        \b11_OFWNT9L_8tZ[46] , \b11_OFWNT9L_8tZ[45] , 
        \b11_OFWNT9L_8tZ[44] , \b11_OFWNT9L_8tZ[43] , 
        \b11_OFWNT9L_8tZ[42] , \b11_OFWNT9L_8tZ[41] , 
        \b11_OFWNT9L_8tZ[40] , \b11_OFWNT9L_8tZ[39] , 
        \b11_OFWNT9L_8tZ[38] , \b11_OFWNT9L_8tZ[37] , 
        \b11_OFWNT9L_8tZ[36] , \b11_OFWNT9L_8tZ[35] , 
        \b11_OFWNT9L_8tZ[34] , \b11_OFWNT9L_8tZ[33] , 
        \b11_OFWNT9L_8tZ[32] , \b11_OFWNT9L_8tZ[31] , 
        \b11_OFWNT9L_8tZ[30] , \b11_OFWNT9L_8tZ[29] , 
        \b11_OFWNT9L_8tZ[28] , \b11_OFWNT9L_8tZ[27] , 
        \b11_OFWNT9L_8tZ[26] , \b11_OFWNT9L_8tZ[25] , 
        \b11_OFWNT9L_8tZ[24] , \b11_OFWNT9L_8tZ[23] , 
        \b11_OFWNT9L_8tZ[22] , \b11_OFWNT9L_8tZ[21] , 
        \b11_OFWNT9L_8tZ[20] , \b11_OFWNT9L_8tZ[19] , 
        \b11_OFWNT9L_8tZ[18] , \b11_OFWNT9L_8tZ[17] , 
        \b11_OFWNT9L_8tZ[16] , \b11_OFWNT9L_8tZ[15] , 
        \b11_OFWNT9L_8tZ[14] , \b11_OFWNT9L_8tZ[13] , 
        \b11_OFWNT9L_8tZ[12] , \b11_OFWNT9L_8tZ[11] , 
        \b11_OFWNT9L_8tZ[10] , \b11_OFWNT9L_8tZ[9] , 
        \b11_OFWNT9L_8tZ[8] , \b11_OFWNT9L_8tZ[7] , 
        \b11_OFWNT9L_8tZ[6] , \b11_OFWNT9L_8tZ[5] , 
        \b11_OFWNT9L_8tZ[4] , \b11_OFWNT9L_8tZ[3] , 
        \b11_OFWNT9L_8tZ[2] , \b11_OFWNT9L_8tZ[1] , 
        \b11_OFWNT9L_8tZ[0] }), .b8_SoWGfWYY(b8_SoWGfWYY), 
        .b8_SoWGfWYY_i(b8_SoWGfWYY_i), .BW_clk_c(BW_clk_c), 
        .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh), .N_44(N_44), 
        .b11_PSyil9s_FMZ(b11_PSyil9s_FMZ), .b4_PLyF(b4_PLyF), 
        .b11_uRrc2XfY_XH(b11_uRrc2XfY_XH), .b13_nUTQBgfDb_Z4D(
        b13_nUTQBgfDb_Z4D), .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), 
        .b16_nYhI39swMeEd_A78(b16_nYhI39swMeEd_A78), 
        .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), .b12_vABZ3qsY_Lyh(
        b12_vABZ3qsY_Lyh), .b11_vABZ3qsY_XH(b11_vABZ3qsY_XH), 
        .b7_PSyi3wy(b7_PSyi3wy), .b8_PSyiBgYG(b8_PSyiBgYG));
    SLE \mdiclink_reg[109]  (.D(temp_count[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[109]_net_1 ));
    SLE \mdiclink_reg[59]  (.D(temp2[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[59]_net_1 ));
    SLE \mdiclink_reg[23]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[23]_net_1 ));
    SLE \mdiclink_reg[6]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[6]_net_1 ));
    SLE \mdiclink_reg[124]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[124]_net_1 ));
    SLE \mdiclink_reg[11]  (.D(freq_14), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[11]_net_1 ));
    SLE \mdiclink_reg[143]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[143]_net_1 ));
    SLE \mdiclink_reg[131]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[131]_net_1 ));
    SLE \mdiclink_reg[9]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[9]_net_1 ));
    SLE \mdiclink_reg[28]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[28]_net_1 ));
    SLE \mdiclink_reg[107]  (.D(temp_count[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[107]_net_1 ));
    SLE \mdiclink_reg[106]  (.D(temp_count[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[106]_net_1 ));
    SLE \mdiclink_reg[100]  (.D(temp_count[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[100]_net_1 ));
    SLE \mdiclink_reg[26]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[26]_net_1 ));
    SLE \mdiclink_reg[71]  (.D(temp3[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[71]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \mdiclink_reg[55]  (.D(temp2[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[55]_net_1 ));
    SLE \mdiclink_reg[13]  (.D(VCC_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[13]_net_1 ));
    SLE \mdiclink_reg[132]  (.D(freq_15), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[132]_net_1 ));
    SLE \mdiclink_reg[62]  (.D(temp2[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[62]_net_1 ));
    SLE \mdiclink_reg[145]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[145]_net_1 ));
    SLE \mdiclink_reg[154]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[154]_net_1 ));
    SLE \mdiclink_reg[18]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[18]_net_1 ));
    SLE \mdiclink_reg[8]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[8]_net_1 ));
    SLE \mdiclink_reg[50]  (.D(temp2[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[50]_net_1 ));
    SLE \mdiclink_reg[73]  (.D(temp3[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[73]_net_1 ));
    SLE \mdiclink_reg[16]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[16]_net_1 ));
    SLE \mdiclink_reg[64]  (.D(temp2[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[64]_net_1 ));
    SLE \mdiclink_reg[57]  (.D(temp2[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[57]_net_1 ));
    SLE \mdiclink_reg[78]  (.D(temp3[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[78]_net_1 ));
    SLE \mdiclink_reg[32]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[32]_net_1 ));
    SLE \mdiclink_reg[149]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[149]_net_1 ));
    SLE \mdiclink_reg[76]  (.D(temp3[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[76]_net_1 ));
    b11_OFWNT9s_8tZ_Z2_x b3_SoW_0 (.b11_OFWNT9L_8tZ({
        \b11_OFWNT9L_8tZ[154] , \b11_OFWNT9L_8tZ[153] , 
        \b11_OFWNT9L_8tZ[152] , \b11_OFWNT9L_8tZ[151] , 
        \b11_OFWNT9L_8tZ[150] , \b11_OFWNT9L_8tZ[149] , 
        \b11_OFWNT9L_8tZ[148] , \b11_OFWNT9L_8tZ[147] , 
        \b11_OFWNT9L_8tZ[146] , \b11_OFWNT9L_8tZ[145] , 
        \b11_OFWNT9L_8tZ[144] , \b11_OFWNT9L_8tZ[143] , 
        \b11_OFWNT9L_8tZ[142] , \b11_OFWNT9L_8tZ[141] , 
        \b11_OFWNT9L_8tZ[140] , \b11_OFWNT9L_8tZ[139] , 
        \b11_OFWNT9L_8tZ[138] , \b11_OFWNT9L_8tZ[137] , 
        \b11_OFWNT9L_8tZ[136] , \b11_OFWNT9L_8tZ[135] , 
        \b11_OFWNT9L_8tZ[134] , \b11_OFWNT9L_8tZ[133] , 
        \b11_OFWNT9L_8tZ[132] , \b11_OFWNT9L_8tZ[131] , 
        \b11_OFWNT9L_8tZ[130] , \b11_OFWNT9L_8tZ[129] , 
        \b11_OFWNT9L_8tZ[128] , \b11_OFWNT9L_8tZ[127] , 
        \b11_OFWNT9L_8tZ[126] , \b11_OFWNT9L_8tZ[125] , 
        \b11_OFWNT9L_8tZ[124] , \b11_OFWNT9L_8tZ[123] , 
        \b11_OFWNT9L_8tZ[122] , \b11_OFWNT9L_8tZ[121] , 
        \b11_OFWNT9L_8tZ[120] , \b11_OFWNT9L_8tZ[119] , 
        \b11_OFWNT9L_8tZ[118] , \b11_OFWNT9L_8tZ[117] , 
        \b11_OFWNT9L_8tZ[116] , \b11_OFWNT9L_8tZ[115] , 
        \b11_OFWNT9L_8tZ[114] , \b11_OFWNT9L_8tZ[113] , 
        \b11_OFWNT9L_8tZ[112] , \b11_OFWNT9L_8tZ[111] , 
        \b11_OFWNT9L_8tZ[110] , \b11_OFWNT9L_8tZ[109] , 
        \b11_OFWNT9L_8tZ[108] , \b11_OFWNT9L_8tZ[107] , 
        \b11_OFWNT9L_8tZ[106] , \b11_OFWNT9L_8tZ[105] , 
        \b11_OFWNT9L_8tZ[104] , \b11_OFWNT9L_8tZ[103] , 
        \b11_OFWNT9L_8tZ[102] , \b11_OFWNT9L_8tZ[101] , 
        \b11_OFWNT9L_8tZ[100] , \b11_OFWNT9L_8tZ[99] , 
        \b11_OFWNT9L_8tZ[98] , \b11_OFWNT9L_8tZ[97] , 
        \b11_OFWNT9L_8tZ[96] , \b11_OFWNT9L_8tZ[95] , 
        \b11_OFWNT9L_8tZ[94] , \b11_OFWNT9L_8tZ[93] , 
        \b11_OFWNT9L_8tZ[92] , \b11_OFWNT9L_8tZ[91] , 
        \b11_OFWNT9L_8tZ[90] , \b11_OFWNT9L_8tZ[89] , 
        \b11_OFWNT9L_8tZ[88] , \b11_OFWNT9L_8tZ[87] , 
        \b11_OFWNT9L_8tZ[86] , \b11_OFWNT9L_8tZ[85] , 
        \b11_OFWNT9L_8tZ[84] , \b11_OFWNT9L_8tZ[83] , 
        \b11_OFWNT9L_8tZ[82] , \b11_OFWNT9L_8tZ[81] , 
        \b11_OFWNT9L_8tZ[80] , \b11_OFWNT9L_8tZ[79] , 
        \b11_OFWNT9L_8tZ[78] , \b11_OFWNT9L_8tZ[77] , 
        \b11_OFWNT9L_8tZ[76] , \b11_OFWNT9L_8tZ[75] , 
        \b11_OFWNT9L_8tZ[74] , \b11_OFWNT9L_8tZ[73] , 
        \b11_OFWNT9L_8tZ[72] , \b11_OFWNT9L_8tZ[71] , 
        \b11_OFWNT9L_8tZ[70] , \b11_OFWNT9L_8tZ[69] , 
        \b11_OFWNT9L_8tZ[68] , \b11_OFWNT9L_8tZ[67] , 
        \b11_OFWNT9L_8tZ[66] , \b11_OFWNT9L_8tZ[65] , 
        \b11_OFWNT9L_8tZ[64] , \b11_OFWNT9L_8tZ[63] , 
        \b11_OFWNT9L_8tZ[62] , \b11_OFWNT9L_8tZ[61] , 
        \b11_OFWNT9L_8tZ[60] , \b11_OFWNT9L_8tZ[59] , 
        \b11_OFWNT9L_8tZ[58] , \b11_OFWNT9L_8tZ[57] , 
        \b11_OFWNT9L_8tZ[56] , \b11_OFWNT9L_8tZ[55] , 
        \b11_OFWNT9L_8tZ[54] , \b11_OFWNT9L_8tZ[53] , 
        \b11_OFWNT9L_8tZ[52] , \b11_OFWNT9L_8tZ[51] , 
        \b11_OFWNT9L_8tZ[50] , \b11_OFWNT9L_8tZ[49] , 
        \b11_OFWNT9L_8tZ[48] , \b11_OFWNT9L_8tZ[47] , 
        \b11_OFWNT9L_8tZ[46] , \b11_OFWNT9L_8tZ[45] , 
        \b11_OFWNT9L_8tZ[44] , \b11_OFWNT9L_8tZ[43] , 
        \b11_OFWNT9L_8tZ[42] , \b11_OFWNT9L_8tZ[41] , 
        \b11_OFWNT9L_8tZ[40] , \b11_OFWNT9L_8tZ[39] , 
        \b11_OFWNT9L_8tZ[38] , \b11_OFWNT9L_8tZ[37] , 
        \b11_OFWNT9L_8tZ[36] , \b11_OFWNT9L_8tZ[35] , 
        \b11_OFWNT9L_8tZ[34] , \b11_OFWNT9L_8tZ[33] , 
        \b11_OFWNT9L_8tZ[32] , \b11_OFWNT9L_8tZ[31] , 
        \b11_OFWNT9L_8tZ[30] , \b11_OFWNT9L_8tZ[29] , 
        \b11_OFWNT9L_8tZ[28] , \b11_OFWNT9L_8tZ[27] , 
        \b11_OFWNT9L_8tZ[26] , \b11_OFWNT9L_8tZ[25] , 
        \b11_OFWNT9L_8tZ[24] , \b11_OFWNT9L_8tZ[23] , 
        \b11_OFWNT9L_8tZ[22] , \b11_OFWNT9L_8tZ[21] , 
        \b11_OFWNT9L_8tZ[20] , \b11_OFWNT9L_8tZ[19] , 
        \b11_OFWNT9L_8tZ[18] , \b11_OFWNT9L_8tZ[17] , 
        \b11_OFWNT9L_8tZ[16] , \b11_OFWNT9L_8tZ[15] , 
        \b11_OFWNT9L_8tZ[14] , \b11_OFWNT9L_8tZ[13] , 
        \b11_OFWNT9L_8tZ[12] , \b11_OFWNT9L_8tZ[11] , 
        \b11_OFWNT9L_8tZ[10] , \b11_OFWNT9L_8tZ[9] , 
        \b11_OFWNT9L_8tZ[8] , \b11_OFWNT9L_8tZ[7] , 
        \b11_OFWNT9L_8tZ[6] , \b11_OFWNT9L_8tZ[5] , 
        \b11_OFWNT9L_8tZ[4] , \b11_OFWNT9L_8tZ[3] , 
        \b11_OFWNT9L_8tZ[2] , \b11_OFWNT9L_8tZ[1] , 
        \b11_OFWNT9L_8tZ[0] }), .mdiclink_reg({
        \mdiclink_reg[154]_net_1 , \mdiclink_reg[153]_net_1 , 
        \mdiclink_reg[152]_net_1 , \mdiclink_reg[151]_net_1 , 
        \mdiclink_reg[150]_net_1 , \mdiclink_reg[149]_net_1 , 
        \mdiclink_reg[148]_net_1 , \mdiclink_reg[147]_net_1 , 
        \mdiclink_reg[146]_net_1 , \mdiclink_reg[145]_net_1 , 
        \mdiclink_reg[144]_net_1 , \mdiclink_reg[143]_net_1 , 
        \mdiclink_reg[142]_net_1 , \mdiclink_reg[141]_net_1 , 
        \mdiclink_reg[140]_net_1 , \mdiclink_reg[139]_net_1 , 
        \mdiclink_reg[138]_net_1 , \mdiclink_reg[137]_net_1 , 
        \mdiclink_reg[136]_net_1 , \mdiclink_reg[135]_net_1 , 
        \mdiclink_reg[134]_net_1 , \mdiclink_reg[133]_net_1 , 
        \mdiclink_reg[132]_net_1 , \mdiclink_reg[131]_net_1 , 
        \mdiclink_reg[130]_net_1 , \mdiclink_reg[129]_net_1 , 
        \mdiclink_reg[128]_net_1 , \mdiclink_reg[127]_net_1 , 
        \mdiclink_reg[126]_net_1 , \mdiclink_reg[125]_net_1 , 
        \mdiclink_reg[124]_net_1 , \mdiclink_reg[123]_net_1 , 
        \mdiclink_reg[122]_net_1 , \mdiclink_reg[121]_net_1 , 
        \mdiclink_reg[120]_net_1 , \mdiclink_reg[119]_net_1 , 
        \mdiclink_reg[118]_net_1 , \mdiclink_reg[117]_net_1 , 
        \mdiclink_reg[116]_net_1 , \mdiclink_reg[115]_net_1 , 
        \mdiclink_reg[114]_net_1 , \mdiclink_reg[113]_net_1 , 
        \mdiclink_reg[112]_net_1 , \mdiclink_reg[111]_net_1 , 
        \mdiclink_reg[110]_net_1 , \mdiclink_reg[109]_net_1 , 
        \mdiclink_reg[108]_net_1 , \mdiclink_reg[107]_net_1 , 
        \mdiclink_reg[106]_net_1 , \mdiclink_reg[105]_net_1 , 
        \mdiclink_reg[104]_net_1 , \mdiclink_reg[103]_net_1 , 
        \mdiclink_reg[102]_net_1 , \mdiclink_reg[101]_net_1 , 
        \mdiclink_reg[100]_net_1 , \mdiclink_reg[99]_net_1 , 
        \mdiclink_reg[98]_net_1 , \mdiclink_reg[97]_net_1 , 
        \mdiclink_reg[96]_net_1 , \mdiclink_reg[95]_net_1 , 
        \mdiclink_reg[94]_net_1 , \mdiclink_reg[93]_net_1 , 
        \mdiclink_reg[92]_net_1 , \mdiclink_reg[91]_net_1 , 
        \mdiclink_reg[90]_net_1 , \mdiclink_reg[89]_net_1 , 
        \mdiclink_reg[88]_net_1 , \mdiclink_reg[87]_net_1 , 
        \mdiclink_reg[86]_net_1 , \mdiclink_reg[85]_net_1 , 
        \mdiclink_reg[84]_net_1 , \mdiclink_reg[83]_net_1 , 
        \mdiclink_reg[82]_net_1 , \mdiclink_reg[81]_net_1 , 
        \mdiclink_reg[80]_net_1 , \mdiclink_reg[79]_net_1 , 
        \mdiclink_reg[78]_net_1 , \mdiclink_reg[77]_net_1 , 
        \mdiclink_reg[76]_net_1 , \mdiclink_reg[75]_net_1 , 
        \mdiclink_reg[74]_net_1 , \mdiclink_reg[73]_net_1 , 
        \mdiclink_reg[72]_net_1 , \mdiclink_reg[71]_net_1 , 
        \mdiclink_reg[70]_net_1 , \mdiclink_reg[69]_net_1 , 
        \mdiclink_reg[68]_net_1 , \mdiclink_reg[67]_net_1 , 
        \mdiclink_reg[66]_net_1 , \mdiclink_reg[65]_net_1 , 
        \mdiclink_reg[64]_net_1 , \mdiclink_reg[63]_net_1 , 
        \mdiclink_reg[62]_net_1 , \mdiclink_reg[61]_net_1 , 
        \mdiclink_reg[60]_net_1 , \mdiclink_reg[59]_net_1 , 
        \mdiclink_reg[58]_net_1 , \mdiclink_reg[57]_net_1 , 
        \mdiclink_reg[56]_net_1 , \mdiclink_reg[55]_net_1 , 
        \mdiclink_reg[54]_net_1 , \mdiclink_reg[53]_net_1 , 
        \mdiclink_reg[52]_net_1 , \mdiclink_reg[51]_net_1 , 
        \mdiclink_reg[50]_net_1 , \mdiclink_reg[49]_net_1 , 
        \mdiclink_reg[48]_net_1 , \mdiclink_reg[47]_net_1 , 
        \mdiclink_reg[46]_net_1 , \mdiclink_reg[45]_net_1 , 
        \mdiclink_reg[44]_net_1 , \mdiclink_reg[43]_net_1 , 
        \mdiclink_reg[42]_net_1 , \mdiclink_reg[41]_net_1 , 
        \mdiclink_reg[40]_net_1 , \mdiclink_reg[39]_net_1 , 
        \mdiclink_reg[38]_net_1 , \mdiclink_reg[37]_net_1 , 
        \mdiclink_reg[36]_net_1 , \mdiclink_reg[35]_net_1 , 
        \mdiclink_reg[34]_net_1 , \mdiclink_reg[33]_net_1 , 
        \mdiclink_reg[32]_net_1 , \mdiclink_reg[31]_net_1 , 
        \mdiclink_reg[30]_net_1 , \mdiclink_reg[29]_net_1 , 
        \mdiclink_reg[28]_net_1 , \mdiclink_reg[27]_net_1 , 
        \mdiclink_reg[26]_net_1 , \mdiclink_reg[25]_net_1 , 
        \mdiclink_reg[24]_net_1 , \mdiclink_reg[23]_net_1 , 
        \mdiclink_reg[22]_net_1 , \mdiclink_reg[21]_net_1 , 
        \mdiclink_reg[20]_net_1 , \mdiclink_reg[19]_net_1 , 
        \mdiclink_reg[18]_net_1 , \mdiclink_reg[17]_net_1 , 
        \mdiclink_reg[16]_net_1 , \mdiclink_reg[15]_net_1 , 
        \mdiclink_reg[14]_net_1 , \mdiclink_reg[13]_net_1 , 
        \mdiclink_reg[12]_net_1 , \mdiclink_reg[11]_net_1 , 
        \mdiclink_reg[10]_net_1 , \mdiclink_reg[9]_net_1 , 
        \mdiclink_reg[8]_net_1 , \mdiclink_reg[7]_net_1 , 
        \mdiclink_reg[6]_net_1 , \mdiclink_reg[5]_net_1 , 
        \mdiclink_reg[4]_net_1 , \mdiclink_reg[3]_net_1 , 
        \mdiclink_reg[2]_net_1 , \mdiclink_reg[1]_net_1 , 
        \mdiclink_reg[0]_net_1 }), .b13_nAzGfFM_sLsv3({
        \b13_nAzGfFM_sLsv3[1] }), .IICE_comm2iice_11(
        IICE_comm2iice[11]), .IICE_comm2iice_0(IICE_comm2iice[0]), 
        .IICE_comm2iice_4(IICE_comm2iice[4]), .IICE_comm2iice_10(
        IICE_comm2iice[10]), .IICE_comm2iice_5(IICE_comm2iice[5]), 
        .IICE_comm2iice_9(IICE_comm2iice[9]), .IICE_comm2iice_1(
        IICE_comm2iice[1]), .IICE_comm2iice_3(IICE_comm2iice[3]), 
        .IICE_comm2iice_2(IICE_comm2iice[2]), .IICE_comm2iice_6(
        IICE_comm2iice[6]), .BW_clk_c(BW_clk_c), .b11_PSyil9s_FMZ(
        b11_PSyil9s_FMZ), .b8_SoWGfWYY_i(b8_SoWGfWYY_i), .b8_SoWGfWYY(
        b8_SoWGfWYY), .b7_yYh03wy(b7_yYh03wy), .b10_OFWNT9khFt(
        b10_OFWNT9khFt), .b9_OFWNT9Mxf(b9_OFWNT9Mxf), .N_44(N_44));
    SLE \mdiclink_reg[91]  (.D(temp_count[24]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[91]_net_1 ));
    SLE \mdiclink_reg[111]  (.D(temp_count[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[111]_net_1 ));
    SLE \mdiclink_reg[147]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[147]_net_1 ));
    SLE \mdiclink_reg[34]  (.D(temp1[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[34]_net_1 ));
    SLE \mdiclink_reg[146]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[146]_net_1 ));
    SLE \mdiclink_reg[140]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[140]_net_1 ));
    b3_uKr_x b8_uKr_IFLY (.b13_nvmFL_fx2rbuQ({IICE_comm2iice[0], 
        IICE_comm2iice[1], IICE_comm2iice[2], IICE_comm2iice[3], 
        IICE_comm2iice[4], IICE_comm2iice[5]}), .b11_uRrc_9urXBb(
        IICE_comm2iice[6]), .b3_PLy(IICE_comm2iice[7]), .b3_PLF(
        IICE_iice2comm), .b7_PLy_PlM(b4_PLyF), .b12_PSyiBgfDb_bd(
        b8_PSyiBgYG), .b12_PSyi2XfYF_bd(b8_PSyi2XYG), 
        .b14_OFWNT9khWqH_3i(b10_OFWNT9khFt), .b13_PSyiBgfDb_Z4D(
        b7_PSyi3wy), .b13_PSyi2XfYF_Z4D(GND_net_1), 
        .b15_OFWNT9khWqH_R9k(b9_OFWNT9Mxf), .b7_yYh03wy(b7_yYh03wy), 
        .b12_nUTQBgfDb_bd(b12_nUTQBgfDb_bd), .b11_uRrc2XfY_XH(
        b11_uRrc2XfY_XH), .b13_nUTQBgfDb_Z4D(b13_nUTQBgfDb_Z4D), 
        .b15_nYhI39swMeEd_Mg(b15_nYhI39swMeEd_Mg), 
        .b16_nYhI39swMeEd_A78(b16_nYhI39swMeEd_A78), .b11_vABZ3qsY_XH(
        b11_vABZ3qsY_XH), .b12_vABZ3qsY_Lyh(b12_vABZ3qsY_Lyh), 
        .b12_ibScJX_E2_bd(b12_ibScJX_E2_bd), .b13_ibScJX_E2_Z4D(
        GND_net_1), .b12_uRrc2XfY_Lyh(b12_uRrc2XfY_Lyh));
    SLE \mdiclink_reg[1]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[1]_net_1 ));
    SLE \mdiclink_reg[93]  (.D(temp_count[22]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[93]_net_1 ));
    SLE \mdiclink_reg[69]  (.D(temp3[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[69]_net_1 ));
    SLE \mdiclink_reg[104]  (.D(temp_count[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[104]_net_1 ));
    SLE \mdiclink_reg[112]  (.D(temp_count[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[112]_net_1 ));
    SLE \mdiclink_reg[22]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[22]_net_1 ));
    SLE \mdiclink_reg[98]  (.D(temp_count[17]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[98]_net_1 ));
    SLE \mdiclink_reg[81]  (.D(temp3[1]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[81]_net_1 ));
    SLE \mdiclink_reg[121]  (.D(temp_sck_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[121]_net_1 ));
    SLE \mdiclink_reg[96]  (.D(temp_count[19]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[96]_net_1 ));
    SLE \mdiclink_reg[138]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[138]_net_1 ));
    SLE \mdiclink_reg[65]  (.D(temp2[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[65]_net_1 ));
    SLE \mdiclink_reg[24]  (.D(freq_1), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[24]_net_1 ));
    SLE \mdiclink_reg[39]  (.D(temp1[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[39]_net_1 ));
    SLE \mdiclink_reg[83]  (.D(temp3_csn_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[83]_net_1 ));
    SLE \mdiclink_reg[12]  (.D(freq_13), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[12]_net_1 ));
    SLE \mdiclink_reg[122]  (.D(temp_so_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[122]_net_1 ));
    SLE \mdiclink_reg[60]  (.D(temp2[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[60]_net_1 ));
    SLE \mdiclink_reg[41]  (.D(temp1[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[41]_net_1 ));
    SLE \mdiclink_reg[151]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[151]_net_1 ));
    SLE \mdiclink_reg[67]  (.D(temp3[15]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[67]_net_1 ));
    SLE \mdiclink_reg[88]  (.D(temp_count[27]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[88]_net_1 ));
    SLE \mdiclink_reg[4]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[4]_net_1 ));
    SLE \mdiclink_reg[72]  (.D(temp3[10]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[72]_net_1 ));
    SLE \mdiclink_reg[86]  (.D(temp_count[29]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[86]_net_1 ));
    SLE \mdiclink_reg[14]  (.D(freq_11), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[14]_net_1 ));
    SLE \mdiclink_reg[35]  (.D(temp1[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[35]_net_1 ));
    SLE \mdiclink_reg[133]  (.D(freq_14), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[133]_net_1 ));
    SLE \mdiclink_reg[43]  (.D(temp1[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[43]_net_1 ));
    SLE \mdiclink_reg[152]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[152]_net_1 ));
    SLE \mdiclink_reg[144]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[144]_net_1 ));
    SLE \mdiclink_reg[74]  (.D(temp3[8]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[74]_net_1 ));
    SLE \mdiclink_reg[29]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[29]_net_1 ));
    SLE \mdiclink_reg[30]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[30]_net_1 ));
    SLE \mdiclink_reg[48]  (.D(temp1[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[48]_net_1 ));
    SLE \mdiclink_reg[37]  (.D(temp1[11]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[37]_net_1 ));
    SLE \mdiclink_reg[46]  (.D(temp1[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[46]_net_1 ));
    SLE \mdiclink_reg[135]  (.D(VCC_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[135]_net_1 ));
    SLE \mdiclink_reg[118]  (.D(temp_count_data[2]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[118]_net_1 ));
    SLE \mdiclink_reg[5]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[5]_net_1 ));
    SLE \mdiclink_reg[19]  (.D(freq_6), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[19]_net_1 ));
    SLE \mdiclink_reg[92]  (.D(temp_count[23]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[92]_net_1 ));
    SLE \mdiclink_reg[25]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[25]_net_1 ));
    SLE \mdiclink_reg[3]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[3]_net_1 ));
    SLE \mdiclink_reg[101]  (.D(temp_count[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[101]_net_1 ));
    SLE \mdiclink_reg[139]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[139]_net_1 ));
    SLE \mdiclink_reg[79]  (.D(temp3[3]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[79]_net_1 ));
    SLE \mdiclink_reg[20]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[20]_net_1 ));
    SLE \mdiclink_reg[94]  (.D(temp_count[21]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[94]_net_1 ));
    SLE \mdiclink_reg[27]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[27]_net_1 ));
    SLE \mdiclink_reg[128]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[128]_net_1 ));
    SLE \mdiclink_reg[51]  (.D(temp2[14]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[51]_net_1 ));
    SLE \mdiclink_reg[15]  (.D(freq_10), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[15]_net_1 ));
    SLE \mdiclink_reg[102]  (.D(temp_count[13]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[102]_net_1 ));
    SLE \mdiclink_reg[113]  (.D(temp_count[2]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[113]_net_1 ));
    SLE \mdiclink_reg[137]  (.D(freq_10), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[137]_net_1 ));
    SLE \mdiclink_reg[136]  (.D(freq_11), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[136]_net_1 ));
    SLE \mdiclink_reg[82]  (.D(temp3[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[82]_net_1 ));
    SLE \mdiclink_reg[130]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[130]_net_1 ));
    SLE \mdiclink_reg[10]  (.D(freq_15), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[10]_net_1 ));
    SLE \mdiclink_reg[75]  (.D(temp3[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[75]_net_1 ));
    SLE \mdiclink_reg[0]  (.D(temp_sck_c), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[0]_net_1 ));
    SLE \mdiclink_reg[53]  (.D(temp2[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[53]_net_1 ));
    SLE \mdiclink_reg[17]  (.D(freq_0), .CLK(BW_clk_c), .EN(VCC_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[17]_net_1 ));
    SLE \mdiclink_reg[115]  (.D(temp_count[0]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[115]_net_1 ));
    SLE \mdiclink_reg[84]  (.D(temp_count[31]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[84]_net_1 ));
    SLE \mdiclink_reg[58]  (.D(temp2[7]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[58]_net_1 ));
    SLE \mdiclink_reg[70]  (.D(temp3[12]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[70]_net_1 ));
    SLE \mdiclink_reg[123]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[123]_net_1 ));
    SLE \mdiclink_reg[77]  (.D(temp3[5]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[77]_net_1 ));
    SLE \mdiclink_reg[56]  (.D(temp2[9]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[56]_net_1 ));
    SLE \mdiclink_reg[99]  (.D(temp_count[16]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[99]_net_1 ));
    SLE \mdiclink_reg[42]  (.D(temp1[6]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[42]_net_1 ));
    SLE \mdiclink_reg[141]  (.D(freq_6), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[141]_net_1 ));
    SLE \mdiclink_reg[7]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[7]_net_1 ));
    SLE \mdiclink_reg[119]  (.D(temp_count_data[1]), .CLK(BW_clk_c), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \mdiclink_reg[119]_net_1 ));
    SLE \mdiclink_reg[44]  (.D(temp1[4]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[44]_net_1 ));
    SLE \mdiclink_reg[125]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[125]_net_1 ));
    SLE \mdiclink_reg[95]  (.D(temp_count[20]), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[95]_net_1 ));
    SLE \mdiclink_reg[153]  (.D(GND_net_1), .CLK(BW_clk_c), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[153]_net_1 ));
    SLE \mdiclink_reg[142]  (.D(freq_2), .CLK(BW_clk_c), .EN(VCC_net_1)
        , .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\mdiclink_reg[142]_net_1 ));
    
endmodule


module b9_ORbIwXaEF_32s_2486674598_0s_x_0(
       b3_ORb_0,
       tck,
       b6_nv_0CC,
       b10_nv_ywKMm9X,
       b12_ORbIwXaEF_bd,
       b8_nv_ZmCtY
    );
output b3_ORb_0;
input  tck;
input  b6_nv_0CC;
input  b10_nv_ywKMm9X;
input  b12_ORbIwXaEF_bd;
input  b8_nv_ZmCtY;

    wire b3_ORb_7_net_1, N_458_i, \b3_ORb[23]_net_1 , VCC_net_1, 
        \b3_ORb[24]_net_1 , \b3_ORb_or[7]_net_1 , GND_net_1, 
        \b3_ORb[25]_net_1 , \b3_ORb[26]_net_1 , \b3_ORb[27]_net_1 , 
        \b3_ORb[28]_net_1 , \b3_ORb[29]_net_1 , \b3_ORb[30]_net_1 , 
        \b3_ORb[31]_net_1 , \b3_ORb[32]_net_1 , \b3_ORb[8]_net_1 , 
        \b3_ORb[9]_net_1 , \b3_ORb[10]_net_1 , \b3_ORb[11]_net_1 , 
        \b3_ORb[12]_net_1 , \b3_ORb[13]_net_1 , \b3_ORb[14]_net_1 , 
        \b3_ORb[15]_net_1 , \b3_ORb[16]_net_1 , \b3_ORb[17]_net_1 , 
        \b3_ORb[18]_net_1 , \b3_ORb[19]_net_1 , \b3_ORb[20]_net_1 , 
        \b3_ORb[21]_net_1 , \b3_ORb[22]_net_1 , \b3_ORb[2]_net_1 , 
        \b3_ORb[3]_net_1 , \b3_ORb[4]_net_1 , \b3_ORb[5]_net_1 , 
        \b3_ORb[6]_net_1 , \b3_ORb[7]_net_1 , un1_b3_ORb9_i_0;
    
    SLE \b3_ORb[7]  (.D(\b3_ORb[8]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[7]_net_1 ));
    SLE \b3_ORb[9]  (.D(\b3_ORb[10]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[9]_net_1 ));
    SLE \b3_ORb[3]  (.D(\b3_ORb[4]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[3]_net_1 ));
    SLE \b3_ORb[23]  (.D(\b3_ORb[24]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[23]_net_1 ));
    SLE \b3_ORb[22]  (.D(\b3_ORb[23]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[22]_net_1 ));
    SLE \b3_ORb[1]  (.D(\b3_ORb[2]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(b3_ORb_0));
    SLE \b3_ORb[10]  (.D(\b3_ORb[11]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[10]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_458_i_0 (.A(b3_ORb_7_net_1), .Y(N_458_i));
    CFG2 #( .INIT(4'hE) )  \b3_ORb_or[7]  (.A(b3_ORb_7_net_1), .B(
        un1_b3_ORb9_i_0), .Y(\b3_ORb_or[7]_net_1 ));
    SLE \b3_ORb[16]  (.D(\b3_ORb[17]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[16]_net_1 ));
    SLE \b3_ORb[11]  (.D(\b3_ORb[12]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[11]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  b3_ORb_7 (.A(b10_nv_ywKMm9X), .B(
        b12_ORbIwXaEF_bd), .Y(b3_ORb_7_net_1));
    SLE \b3_ORb[17]  (.D(\b3_ORb[18]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[17]_net_1 ));
    SLE \b3_ORb[5]  (.D(\b3_ORb[6]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[5]_net_1 ));
    SLE \b3_ORb[28]  (.D(\b3_ORb[29]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[28]_net_1 ));
    SLE \b3_ORb[6]  (.D(\b3_ORb[7]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[6]_net_1 ));
    SLE \b3_ORb[29]  (.D(\b3_ORb[30]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[29]_net_1 ));
    SLE \b3_ORb[13]  (.D(\b3_ORb[14]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[13]_net_1 ));
    SLE \b3_ORb[12]  (.D(\b3_ORb[13]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[12]_net_1 ));
    SLE \b3_ORb[24]  (.D(\b3_ORb[25]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[24]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hC8) )  un1_b3_ORb9_i (.A(b10_nv_ywKMm9X), .B(
        b12_ORbIwXaEF_bd), .C(b8_nv_ZmCtY), .Y(un1_b3_ORb9_i_0));
    SLE \b3_ORb[2]  (.D(\b3_ORb[3]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[2]_net_1 ));
    SLE \b3_ORb[25]  (.D(\b3_ORb[26]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[25]_net_1 ));
    SLE \b3_ORb[30]  (.D(\b3_ORb[31]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[30]_net_1 ));
    SLE \b3_ORb[18]  (.D(\b3_ORb[19]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[18]_net_1 ));
    SLE \b3_ORb[20]  (.D(\b3_ORb[21]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[20]_net_1 ));
    SLE \b3_ORb[19]  (.D(\b3_ORb[20]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[19]_net_1 ));
    SLE \b3_ORb[31]  (.D(\b3_ORb[32]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[31]_net_1 ));
    SLE \b3_ORb[14]  (.D(\b3_ORb[15]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[14]_net_1 ));
    SLE \b3_ORb[26]  (.D(\b3_ORb[27]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[26]_net_1 ));
    SLE \b3_ORb[4]  (.D(\b3_ORb[5]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[4]_net_1 ));
    SLE \b3_ORb[21]  (.D(\b3_ORb[22]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[21]_net_1 ));
    SLE \b3_ORb[8]  (.D(\b3_ORb[9]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[8]_net_1 ));
    SLE \b3_ORb[15]  (.D(\b3_ORb[16]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[15]_net_1 ));
    SLE \b3_ORb[27]  (.D(\b3_ORb[28]_net_1 ), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[27]_net_1 ));
    SLE \b3_ORb[32]  (.D(b6_nv_0CC), .CLK(tck), .EN(
        \b3_ORb_or[7]_net_1 ), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        N_458_i), .SD(VCC_net_1), .LAT(GND_net_1), .Q(
        \b3_ORb[32]_net_1 ));
    
endmodule


module jtag_interface_x_0(
       b11_uRrc_WYOFjZ,
       b11_uRrc_9urXBb,
       dr2_tck_i,
       b9_96_cLqgOF4,
       b10_8Kz_fFfsjX,
       b5_OvyH3,
       b8_nv_ZmCtY,
       b7_nFG0rDY,
       b10_nv_ywKMm9X,
       b6_PLF_Bq,
       hcr_update,
       ch_update,
       b6_nv_0CC,
       atrstb,
       atdo,
       atdi,
       atms,
       atck
    );
input  [0:0] b11_uRrc_WYOFjZ;
output [0:0] b11_uRrc_9urXBb;
output dr2_tck_i;
output b9_96_cLqgOF4;
output b10_8Kz_fFfsjX;
output b5_OvyH3;
output b8_nv_ZmCtY;
output b7_nFG0rDY;
output b10_nv_ywKMm9X;
input  b6_PLF_Bq;
output hcr_update;
output ch_update;
output b6_nv_0CC;
input  atrstb;
output atdo;
input  atdi;
input  atms;
input  atck;

    wire identify_clk_int, \b6_uS_MrX[2] , \b6_uS_MrX[3] , 
        b9_96_cLqgOF4_2, \b6_uS_MrX[0] , \b6_uS_MrX[4] , 
        \b6_uS_MrX[1] , b9_96_cLqgOF3_net_1, b3_1Um, 
        identify_clk2_no_clk_buffer_needed, b9_PLF_6lNa2_net_1, 
        \UIREGdummy[0] , \UIREGdummy[7] , URSTBdummy, GND_net_1, 
        VCC_net_1;
    
    CFG4 #( .INIT(16'h0008) )  b9_96_cLqgOF3 (.A(\b6_uS_MrX[0] ), .B(
        b9_96_cLqgOF4_2), .C(\b6_uS_MrX[4] ), .D(\b6_uS_MrX[1] ), .Y(
        b9_96_cLqgOF3_net_1));
    CFG2 #( .INIT(4'h8) )  b10_8Kz_fFfsjX_inst_1 (.A(b9_96_cLqgOF4), 
        .B(b3_1Um), .Y(b10_8Kz_fFfsjX));
    CFG3 #( .INIT(8'h80) )  b10_nv_ywKMm9X_inst_1 (.A(b3_1Um), .B(
        b9_96_cLqgOF3_net_1), .C(b7_nFG0rDY), .Y(b10_nv_ywKMm9X));
    GND GND (.Y(GND_net_1));
    UJTAG b9_Rcmi_KsDw (.UDRCAP(b7_nFG0rDY), .UDRSH(b5_OvyH3), .UDRUPD(
        identify_clk2_no_clk_buffer_needed), .UIREG({\UIREGdummy[7] , 
        b3_1Um, \b6_uS_MrX[4] , \b6_uS_MrX[3] , \b6_uS_MrX[2] , 
        \b6_uS_MrX[1] , \b6_uS_MrX[0] , \UIREGdummy[0] }), .URSTB(
        URSTBdummy), .UDRCK(identify_clk_int), .UTDI(b6_nv_0CC), .UTDO(
        b9_PLF_6lNa2_net_1), .TDI(atdi), .TMS(atms), .TCK(atck), 
        .TRSTB(atrstb), .TDO(atdo));
    CFG3 #( .INIT(8'h80) )  b8_nv_ZmCtY_inst_1 (.A(b3_1Um), .B(
        b9_96_cLqgOF3_net_1), .C(b5_OvyH3), .Y(b8_nv_ZmCtY));
    CFG3 #( .INIT(8'h80) )  b9_nv_oQwfYF_3 (.A(
        identify_clk2_no_clk_buffer_needed), .B(b9_96_cLqgOF3_net_1), 
        .C(b3_1Um), .Y(ch_update));
    CFG2 #( .INIT(4'h8) )  b10_8Kz_rKlrtX_3 (.A(b10_8Kz_fFfsjX), .B(
        identify_clk2_no_clk_buffer_needed), .Y(hcr_update));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h1) )  b9_96_cLqgOF3_2 (.A(\b6_uS_MrX[2] ), .B(
        \b6_uS_MrX[3] ), .Y(b9_96_cLqgOF4_2));
    CLKINT jtag_clkint_prim (.A(identify_clk_int), .Y(dr2_tck_i));
    CFG4 #( .INIT(16'h0400) )  b9_96_cLqgOF4_inst_1 (.A(\b6_uS_MrX[0] )
        , .B(b9_96_cLqgOF4_2), .C(\b6_uS_MrX[4] ), .D(\b6_uS_MrX[1] ), 
        .Y(b9_96_cLqgOF4));
    CFG3 #( .INIT(8'h80) )  \b11_uRrc_9urXBb[0]  (.A(
        b11_uRrc_WYOFjZ[0]), .B(b3_1Um), .C(b9_96_cLqgOF3_net_1), .Y(
        b11_uRrc_9urXBb[0]));
    CFG4 #( .INIT(16'hC080) )  b9_PLF_6lNa2 (.A(b9_96_cLqgOF4), .B(
        b3_1Um), .C(b6_PLF_Bq), .D(b9_96_cLqgOF3_net_1), .Y(
        b9_PLF_6lNa2_net_1));
    
endmodule


module b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0(
       b11_uRrc_WYOFjZ,
       b13_nvmFL_fx2rbuQ,
       dr2_tck,
       b6_nv_0CC,
       hcr_update,
       b10_8Kz_fFfsjX,
       b12_ORbIwXaEF_bd,
       b9_96_cLqgOF4,
       tdo_sig,
       b7_nFG0rDY,
       b5_OvyH3,
       IICE_iice2comm,
       b6_PLF_Bq
    );
output [0:0] b11_uRrc_WYOFjZ;
output [5:0] b13_nvmFL_fx2rbuQ;
input  dr2_tck;
input  b6_nv_0CC;
input  hcr_update;
input  b10_8Kz_fFfsjX;
output b12_ORbIwXaEF_bd;
input  b9_96_cLqgOF4;
input  tdo_sig;
input  b7_nFG0rDY;
input  b5_OvyH3;
input  IICE_iice2comm;
output b6_PLF_Bq;

    wire \b9_OvyH3_saL[1]_net_1 , VCC_net_1, \b9_OvyH3_saL[2]_net_1 , 
        b9_OvyH3_saL_0_sqmuxa_net_1, GND_net_1, 
        \b9_OvyH3_saL[3]_net_1 , \b9_OvyH3_saL[4]_net_1 , 
        \b9_OvyH3_saL[5]_net_1 , \b9_OvyH3_saL[6]_net_1 , 
        \b9_OvyH3_saL[7]_net_1 , \b9_OvyH3_saL[0]_net_1 , 
        b3_PLF_d_net_1;
    
    SLE \genblk1.b10_dZst39_EF3[5]  (.D(\b9_OvyH3_saL[5]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[4]));
    SLE \genblk1.b10_dZst39_EF3[4]  (.D(\b9_OvyH3_saL[4]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[3]));
    SLE \genblk1.b10_dZst39_EF3[3]  (.D(\b9_OvyH3_saL[3]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[2]));
    SLE \genblk1.b10_dZst39_EF3[1]  (.D(\b9_OvyH3_saL[1]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[0]));
    SLE \b9_OvyH3_saL[6]  (.D(\b9_OvyH3_saL[7]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[6]_net_1 ));
    SLE \b9_OvyH3_saL[3]  (.D(\b9_OvyH3_saL[4]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[3]_net_1 ));
    SLE \genblk1.b10_dZst39_EF3[0]  (.D(\b9_OvyH3_saL[0]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b11_uRrc_WYOFjZ[0]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hFE10) )  b3_PLF (.A(b9_96_cLqgOF4), .B(
        b12_ORbIwXaEF_bd), .C(IICE_iice2comm), .D(b3_PLF_d_net_1), .Y(
        b6_PLF_Bq));
    SLE \genblk1.b10_dZst39_EF3[7]  (.D(\b9_OvyH3_saL[7]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b12_ORbIwXaEF_bd));
    SLE \b9_OvyH3_saL[5]  (.D(\b9_OvyH3_saL[6]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[5]_net_1 ));
    SLE \genblk1.b10_dZst39_EF3[6]  (.D(\b9_OvyH3_saL[6]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[5]));
    SLE \genblk1.b10_dZst39_EF3[2]  (.D(\b9_OvyH3_saL[2]_net_1 ), .CLK(
        hcr_update), .EN(b10_8Kz_fFfsjX), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(b13_nvmFL_fx2rbuQ[1]));
    SLE \b9_OvyH3_saL[7]  (.D(b6_nv_0CC), .CLK(dr2_tck), .EN(
        b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \b9_OvyH3_saL[7]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \b9_OvyH3_saL[1]  (.D(\b9_OvyH3_saL[2]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[1]_net_1 ));
    SLE \b9_OvyH3_saL[0]  (.D(\b9_OvyH3_saL[1]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[0]_net_1 ));
    SLE \b9_OvyH3_saL[4]  (.D(\b9_OvyH3_saL[5]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[4]_net_1 ));
    SLE \b9_OvyH3_saL[2]  (.D(\b9_OvyH3_saL[3]_net_1 ), .CLK(dr2_tck), 
        .EN(b9_OvyH3_saL_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\b9_OvyH3_saL[2]_net_1 ));
    CFG3 #( .INIT(8'h40) )  b9_OvyH3_saL_0_sqmuxa (.A(b7_nFG0rDY), .B(
        b5_OvyH3), .C(b10_8Kz_fFfsjX), .Y(b9_OvyH3_saL_0_sqmuxa_net_1));
    CFG3 #( .INIT(8'hD8) )  b3_PLF_d (.A(b9_96_cLqgOF4), .B(
        \b9_OvyH3_saL[0]_net_1 ), .C(tdo_sig), .Y(b3_PLF_d_net_1));
    
endmodule


module comm_block_x(
       IICE_comm2iice,
       IICE_iice2comm,
       atck,
       atdi,
       atdo,
       atms,
       atrstb
    );
output [0:11] IICE_comm2iice;
input  IICE_iice2comm;
input  atck;
input  atdi;
output atdo;
input  atms;
input  atrstb;

    wire hcr_update, b10_8Kz_fFfsjX, \b11_uRrc_WYOFjZ[0] , 
        b12_ORbIwXaEF_bd, tdo_sig, \jtagi.b7_nFG0rDY , 
        \jtagi.b5_OvyH3 , GND_net_1, VCC_net_1, \jtagi.b9_96_cLqgOF4 , 
        b6_PLF_Bq;
    
    VCC VCC (.Y(VCC_net_1));
    b9_ORbIwXaEF_32s_2486674598_0s_x_0 b9_ORb_xNywD (.b3_ORb_0(tdo_sig)
        , .tck(IICE_comm2iice[11]), .b6_nv_0CC(IICE_comm2iice[7]), 
        .b10_nv_ywKMm9X(IICE_comm2iice[9]), .b12_ORbIwXaEF_bd(
        b12_ORbIwXaEF_bd), .b8_nv_ZmCtY(IICE_comm2iice[10]));
    jtag_interface_x_0 jtagi (.b11_uRrc_WYOFjZ({\b11_uRrc_WYOFjZ[0] }), 
        .b11_uRrc_9urXBb({IICE_comm2iice[6]}), .dr2_tck_i(
        IICE_comm2iice[11]), .b9_96_cLqgOF4(\jtagi.b9_96_cLqgOF4 ), 
        .b10_8Kz_fFfsjX(b10_8Kz_fFfsjX), .b5_OvyH3(\jtagi.b5_OvyH3 ), 
        .b8_nv_ZmCtY(IICE_comm2iice[10]), .b7_nFG0rDY(
        \jtagi.b7_nFG0rDY ), .b10_nv_ywKMm9X(IICE_comm2iice[9]), 
        .b6_PLF_Bq(b6_PLF_Bq), .hcr_update(hcr_update), .ch_update(
        IICE_comm2iice[8]), .b6_nv_0CC(IICE_comm2iice[7]), .atrstb(
        atrstb), .atdo(atdo), .atdi(atdi), .atms(atms), .atck(atck));
    GND GND (.Y(GND_net_1));
    b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0 b7_Rcmi_ql 
        (.b11_uRrc_WYOFjZ({\b11_uRrc_WYOFjZ[0] }), .b13_nvmFL_fx2rbuQ({
        IICE_comm2iice[0], IICE_comm2iice[1], IICE_comm2iice[2], 
        IICE_comm2iice[3], IICE_comm2iice[4], IICE_comm2iice[5]}), 
        .dr2_tck(IICE_comm2iice[11]), .b6_nv_0CC(IICE_comm2iice[7]), 
        .hcr_update(hcr_update), .b10_8Kz_fFfsjX(b10_8Kz_fFfsjX), 
        .b12_ORbIwXaEF_bd(b12_ORbIwXaEF_bd), .b9_96_cLqgOF4(
        \jtagi.b9_96_cLqgOF4 ), .tdo_sig(tdo_sig), .b7_nFG0rDY(
        \jtagi.b7_nFG0rDY ), .b5_OvyH3(\jtagi.b5_OvyH3 ), 
        .IICE_iice2comm(IICE_iice2comm), .b6_PLF_Bq(b6_PLF_Bq));
    
endmodule


module syn_identify_core0_0(
       temp1,
       temp2,
       temp3,
       temp_count_data,
       temp_count,
       freq_1,
       freq_2,
       freq_0,
       freq_6,
       freq_10,
       freq_11,
       freq_13,
       freq_14,
       freq_15,
       atck,
       atdi,
       atdo,
       atms,
       atrstb,
       BW_clk_c,
       temp_sck_c,
       temp1_csn_c,
       temp2_csn_c,
       temp3_csn_c,
       temp_so_c
    );
input  [15:0] temp1;
input  [15:0] temp2;
input  [15:0] temp3;
input  [4:0] temp_count_data;
input  [31:0] temp_count;
input  freq_1;
input  freq_2;
input  freq_0;
input  freq_6;
input  freq_10;
input  freq_11;
input  freq_13;
input  freq_14;
input  freq_15;
input  atck;
input  atdi;
output atdo;
input  atms;
input  atrstb;
input  BW_clk_c;
input  temp_sck_c;
input  temp1_csn_c;
input  temp2_csn_c;
input  temp3_csn_c;
input  temp_so_c;

    wire \IICE_comm2iice[11] , \IICE_comm2iice[10] , 
        \IICE_comm2iice[9] , \IICE_comm2iice[8] , \IICE_comm2iice[7] , 
        \IICE_comm2iice[6] , \IICE_comm2iice[5] , \IICE_comm2iice[4] , 
        \IICE_comm2iice[3] , \IICE_comm2iice[2] , \IICE_comm2iice[1] , 
        \IICE_comm2iice[0] , IICE_iice2comm, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    IICE_x IICE_INST (.temp1({temp1[15], temp1[14], temp1[13], 
        temp1[12], temp1[11], temp1[10], temp1[9], temp1[8], temp1[7], 
        temp1[6], temp1[5], temp1[4], temp1[3], temp1[2], temp1[1], 
        temp1[0]}), .temp2({temp2[15], temp2[14], temp2[13], temp2[12], 
        temp2[11], temp2[10], temp2[9], temp2[8], temp2[7], temp2[6], 
        temp2[5], temp2[4], temp2[3], temp2[2], temp2[1], temp2[0]}), 
        .temp3({temp3[15], temp3[14], temp3[13], temp3[12], temp3[11], 
        temp3[10], temp3[9], temp3[8], temp3[7], temp3[6], temp3[5], 
        temp3[4], temp3[3], temp3[2], temp3[1], temp3[0]}), 
        .temp_count_data({temp_count_data[4], temp_count_data[3], 
        temp_count_data[2], temp_count_data[1], temp_count_data[0]}), 
        .temp_count({temp_count[31], temp_count[30], temp_count[29], 
        temp_count[28], temp_count[27], temp_count[26], temp_count[25], 
        temp_count[24], temp_count[23], temp_count[22], temp_count[21], 
        temp_count[20], temp_count[19], temp_count[18], temp_count[17], 
        temp_count[16], temp_count[15], temp_count[14], temp_count[13], 
        temp_count[12], temp_count[11], temp_count[10], temp_count[9], 
        temp_count[8], temp_count[7], temp_count[6], temp_count[5], 
        temp_count[4], temp_count[3], temp_count[2], temp_count[1], 
        temp_count[0]}), .IICE_comm2iice({\IICE_comm2iice[11] , 
        \IICE_comm2iice[10] , \IICE_comm2iice[9] , \IICE_comm2iice[8] , 
        \IICE_comm2iice[7] , \IICE_comm2iice[6] , \IICE_comm2iice[5] , 
        \IICE_comm2iice[4] , \IICE_comm2iice[3] , \IICE_comm2iice[2] , 
        \IICE_comm2iice[1] , \IICE_comm2iice[0] }), .freq_1(freq_1), 
        .freq_2(freq_2), .freq_0(freq_0), .freq_6(freq_6), .freq_10(
        freq_10), .freq_11(freq_11), .freq_13(freq_13), .freq_14(
        freq_14), .freq_15(freq_15), .BW_clk_c(BW_clk_c), .temp_sck_c(
        temp_sck_c), .temp1_csn_c(temp1_csn_c), .temp2_csn_c(
        temp2_csn_c), .temp3_csn_c(temp3_csn_c), .temp_so_c(temp_so_c), 
        .IICE_iice2comm(IICE_iice2comm));
    GND GND (.Y(GND_net_1));
    comm_block_x comm_block_INST (.IICE_comm2iice({\IICE_comm2iice[0] , 
        \IICE_comm2iice[1] , \IICE_comm2iice[2] , \IICE_comm2iice[3] , 
        \IICE_comm2iice[4] , \IICE_comm2iice[5] , \IICE_comm2iice[6] , 
        \IICE_comm2iice[7] , \IICE_comm2iice[8] , \IICE_comm2iice[9] , 
        \IICE_comm2iice[10] , \IICE_comm2iice[11] }), .IICE_iice2comm(
        IICE_iice2comm), .atck(atck), .atdi(atdi), .atdo(atdo), .atms(
        atms), .atrstb(atrstb));
    
endmodule


module build_sb_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module build_sb_CCC_0_FCCC(
       temp_sck_c,
       temp_sck_c_i_0,
       BW_clk_c,
       BW_clk_c_i_0,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output temp_sck_c;
output temp_sck_c_i_0;
output BW_clk_c;
output BW_clk_c_i_0;
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL2_net, GL1_net, VCC_net_1, GND_net_1;
    
    CLKINT GL1_INST (.A(GL1_net), .Y(temp_sck_c));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  GL1_INST_RNI8343 (.A(temp_sck_c), .Y(
        temp_sck_c_i_0));
    GND GND (.Y(GND_net_1));
    CLKINT GL2_INST (.A(GL2_net), .Y(BW_clk_c));
    CCC #( .INIT(210'h0000007FB8000044564003F0BC2B09C20E739DEFFC4C980C00B01)
        , .VCOFREQUENCY(600.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(), 
        .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(VCC_net_1), 
        .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), .NGMUX1_SEL(
        GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(GND_net_1), 
        .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(VCC_net_1), 
        .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(VCC_net_1), 
        .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(VCC_net_1), 
        .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(VCC_net_1), 
        .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(), .GL1(GL1_net), .GL2(
        GL2_net), .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    CFG1 #( .INIT(2'h1) )  GL2_INST_RNI98ED (.A(BW_clk_c), .Y(
        BW_clk_c_i_0));
    
endmodule


module build_sb(
       temp_sck_c,
       temp_sck_c_i_0,
       BW_clk_c,
       BW_clk_c_i_0
    );
output temp_sck_c;
output temp_sck_c_i_0;
output BW_clk_c;
output BW_clk_c_i_0;

    wire FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, GND_net_1, 
        VCC_net_1;
    
    build_sb_FABOSC_0_OSC FABOSC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    build_sb_CCC_0_FCCC CCC_0 (.temp_sck_c(temp_sck_c), 
        .temp_sck_c_i_0(temp_sck_c_i_0), .BW_clk_c(BW_clk_c), 
        .BW_clk_c_i_0(BW_clk_c_i_0), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    GND GND (.Y(GND_net_1));
    
endmodule


module build(
       BW,
       SENSE_DIN,
       adc_d0,
       BW_out,
       SENSE_DOUT,
       dac1_db,
       fl_a,
       fl_dq,
       ANTF_n1,
       ANTF_n2,
       DEVRST_N,
       GPIO10,
       GPIO11,
       GPIO8,
       GPIO9,
       GPS1_I0,
       GPS1_I1,
       GPS1_LD,
       GPS1_Q0,
       GPS1_Q1,
       GPS2_LD,
       GPS2_Q0,
       GPS2_Q1,
       GPS_I0,
       GPS_I1,
       adc_clk,
       adc_oen,
       adc_of,
       osc_vcc,
       temp_so,
       AMP_EN,
       BW_36,
       BW_clk,
       CSN_n1,
       CTR1,
       CTR2,
       CTR3,
       CTR4,
       CTR5,
       CTR6,
       CTR7,
       GPIO1,
       GPIO12,
       GPIO14,
       GPIO15,
       GPIO16,
       GPIO17,
       GPIO19,
       GPIO2,
       GPIO20,
       GPIO3,
       GPIO4,
       GPIO5,
       GPIO6,
       GPIO7,
       GPS1_IDLE,
       GPS1_PGM,
       GPS1_SCLK,
       GPS1_SDATA,
       GPS1_SHDN,
       REF_CE,
       REF_CLK,
       REF_DATA,
       REF_LD,
       REF_LE,
       REF_MXOUT,
       SENSE_CS_1,
       adc_shdn,
       clk_out_n1,
       clk_out_n2,
       dac1_clk,
       dac1_sleep,
       dac2_clk,
       dsa_clk,
       dsa_data,
       dsa_le,
       en_modul,
       fl_byten,
       fl_cen,
       fl_oen,
       fl_resetn,
       fl_ryby,
       fl_wen,
       fl_wpn,
       oclk_1,
       out1,
       out2,
       sr_cs1n,
       sr_cs2,
       sr_lbn,
       sr_oen,
       sr_ubn,
       sr_wen,
       temp1_csn,
       temp2_csn,
       temp3_csn,
       temp_sck,
       atck,
       atdi,
       atdo,
       atms,
       atrstb
    );
input  [14:0] BW;
input  [1:0] SENSE_DIN;
input  [13:0] adc_d0;
output [14:0] BW_out;
output [1:0] SENSE_DOUT;
output [13:5] dac1_db;
output [25:0] fl_a;
output [7:0] fl_dq;
input  ANTF_n1;
input  ANTF_n2;
input  DEVRST_N;
input  GPIO10;
input  GPIO11;
input  GPIO8;
input  GPIO9;
input  GPS1_I0;
input  GPS1_I1;
input  GPS1_LD;
input  GPS1_Q0;
input  GPS1_Q1;
input  GPS2_LD;
input  GPS2_Q0;
input  GPS2_Q1;
input  GPS_I0;
input  GPS_I1;
input  adc_clk;
input  adc_oen;
input  adc_of;
input  osc_vcc;
input  temp_so;
output AMP_EN;
output BW_36;
output BW_clk;
output CSN_n1;
output CTR1;
output CTR2;
output CTR3;
output CTR4;
output CTR5;
output CTR6;
output CTR7;
output GPIO1;
output GPIO12;
output GPIO14;
output GPIO15;
output GPIO16;
output GPIO17;
output GPIO19;
output GPIO2;
output GPIO20;
output GPIO3;
output GPIO4;
output GPIO5;
output GPIO6;
output GPIO7;
output GPS1_IDLE;
output GPS1_PGM;
output GPS1_SCLK;
output GPS1_SDATA;
output GPS1_SHDN;
output REF_CE;
output REF_CLK;
output REF_DATA;
output REF_LD;
output REF_LE;
output REF_MXOUT;
output SENSE_CS_1;
output adc_shdn;
output clk_out_n1;
output clk_out_n2;
output dac1_clk;
output dac1_sleep;
output dac2_clk;
output dsa_clk;
output dsa_data;
output dsa_le;
output en_modul;
output fl_byten;
output fl_cen;
output fl_oen;
output fl_resetn;
output fl_ryby;
output fl_wen;
output fl_wpn;
output oclk_1;
output out1;
output out2;
output sr_cs1n;
output sr_cs2;
output sr_lbn;
output sr_oen;
output sr_ubn;
output sr_wen;
output temp1_csn;
output temp2_csn;
output temp3_csn;
output temp_sck;
input  atck;
input  atdi;
output atdo;
input  atms;
input  atrstb;

    wire VCC_net_1, GND_net_1, \freq[7] , \freq[8] , \freq[9] , 
        \freq[13] , \freq[17] , \freq[18] , \freq[20] , \freq[21] , 
        \freq[22] , \temp_count_data[0] , \temp_count_data[1] , 
        \temp_count_data[2] , \temp_count_data[3] , 
        \temp_count_data[4] , \temp_count[0] , \temp_count[1] , 
        \temp_count[2] , \temp_count[3] , \temp_count[4] , 
        \temp_count[5] , \temp_count[6] , \temp_count[7] , 
        \temp_count[8] , \temp_count[9] , \temp_count[10] , 
        \temp_count[11] , \temp_count[12] , \temp_count[13] , 
        \temp_count[14] , \temp_count[15] , \temp_count[16] , 
        \temp_count[17] , \temp_count[18] , \temp_count[20] , 
        \temp_count[21] , \temp_count[22] , \temp_count[23] , 
        \temp_count[24] , \temp_count[25] , \temp_count[26] , 
        \temp_count[27] , \temp_count[28] , \temp_count[29] , 
        \temp_count[30] , \temp_count[31] , \temp3[0] , \temp3[1] , 
        \temp3[2] , \temp3[3] , \temp3[4] , \temp3[5] , \temp3[6] , 
        \temp3[7] , \temp3[8] , \temp3[9] , \temp3[10] , \temp3[11] , 
        \temp3[12] , \temp3[13] , \temp3[14] , \temp3[15] , \temp2[0] , 
        \temp2[1] , \temp2[2] , \temp2[3] , \temp2[4] , \temp2[5] , 
        \temp2[6] , \temp2[7] , \temp2[8] , \temp2[9] , \temp2[10] , 
        \temp2[11] , \temp2[12] , \temp2[13] , \temp2[14] , 
        \temp2[15] , \temp1[0] , \temp1[1] , \temp1[2] , \temp1[3] , 
        \temp1[4] , \temp1[5] , \temp1[6] , \temp1[7] , \temp1[8] , 
        \temp1[9] , \temp1[10] , \temp1[11] , \temp1[12] , \temp1[13] , 
        \temp1[14] , \temp1[15] , ANTF_n1_c, ANTF_n2_c, \BW_c[0] , 
        \BW_c[1] , \BW_c[2] , \BW_c[3] , \BW_c[4] , \BW_c[5] , 
        \BW_c[6] , \BW_c[7] , \BW_c[8] , \BW_c[9] , \BW_c[10] , 
        \BW_c[11] , \BW_c[12] , \BW_c[13] , \BW_c[14] , GPIO10_c, 
        GPIO11_c, GPIO8_c, GPIO9_c, GPS1_I0_c, GPS1_I1_c, GPS1_LD_c, 
        GPS1_Q0_c, GPS1_Q1_c, GPS2_LD_c, GPS2_Q0_c, GPS2_Q1_c, 
        GPS_I0_c, GPS_I1_c, GPIO6_c, GPIO4_c, adc_clk_c, \adc_d0_c[0] , 
        \adc_d0_c[1] , \adc_d0_c[2] , \adc_d0_c[3] , \adc_d0_c[4] , 
        \adc_d0_c[5] , \adc_d0_c[6] , \adc_d0_c[7] , \adc_d0_c[8] , 
        \adc_d0_c[9] , \adc_d0_c[10] , \adc_d0_c[11] , \adc_d0_c[12] , 
        \adc_d0_c[13] , adc_oen_c, adc_of_c, osc_vcc_c, temp_so_c, 
        BW_clk_c, \BW_out_c[0] , \BW_out_c[1] , \BW_out_c[2] , 
        \BW_out_c[3] , \BW_out_c[4] , \BW_out_c[5] , \BW_out_c[6] , 
        \BW_out_c[7] , \BW_out_c[8] , \BW_out_c[9] , \BW_out_c[10] , 
        \BW_out_c[11] , \BW_out_c[12] , \BW_out_c[13] , \BW_out_c[14] , 
        GPIO14_c, GPIO16_c, GPIO20_c, GPIO3_c, GPIO5_c, GPIO7_c, 
        SENSE_CS_1_c, \SENSE_DOUT_c[1] , dac1_clk_c, \dac1_db_c[5] , 
        \dac1_db_c[6] , \dac1_db_c[7] , \dac1_db_c[8] , \dac1_db_c[9] , 
        \dac1_db_c[10] , \dac1_db_c[11] , \dac1_db_c[12] , 
        \dac1_db_c[13] , dac2_clk_c, oclk_1_c, temp1_csn_c, 
        temp2_csn_c, temp3_csn_c, temp_sck_c, temp_sck_c_i_0, 
        BW_clk_c_i_0, GPIO9_c_i_0, GPIO8_c_i_0, \temp_count[19] ;
    
    INBUF \BW_ibuf[9]  (.PAD(BW[9]), .Y(\BW_c[9] ));
    INBUF GPS1_I1_ibuf (.PAD(GPS1_I1), .Y(GPS1_I1_c));
    INBUF \BW_ibuf[3]  (.PAD(BW[3]), .Y(\BW_c[3] ));
    INBUF \adc_d0_ibuf[8]  (.PAD(adc_d0[8]), .Y(\adc_d0_c[8] ));
    TRIBUFF \fl_dq_obuft[1]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[1]));
    OUTBUF \BW_out_obuf[7]  (.D(\BW_out_c[7] ), .PAD(BW_out[7]));
    OUTBUF GPIO3_obuf (.D(GPIO3_c), .PAD(GPIO3));
    INBUF \adc_d0_ibuf[6]  (.PAD(adc_d0[6]), .Y(\adc_d0_c[6] ));
    INBUF \BW_ibuf[5]  (.PAD(BW[5]), .Y(\BW_c[5] ));
    OUTBUF \BW_out_obuf[8]  (.D(\BW_out_c[8] ), .PAD(BW_out[8]));
    INBUF GPS2_Q1_ibuf (.PAD(GPS2_Q1), .Y(GPS2_Q1_c));
    led_igloo led_igloo_0 (.temp_count_data({\temp_count_data[4] , 
        \temp_count_data[3] , \temp_count_data[2] , 
        \temp_count_data[1] , \temp_count_data[0] }), .BW_out_c({
        \BW_out_c[14] , \BW_out_c[13] , \BW_out_c[12] , \BW_out_c[11] , 
        \BW_out_c[10] , \BW_out_c[9] , \BW_out_c[8] , \BW_out_c[7] , 
        \BW_out_c[6] , \BW_out_c[5] , \BW_out_c[4] , \BW_out_c[3] , 
        \BW_out_c[2] , \BW_out_c[1] , \BW_out_c[0] }), .BW_c({
        \BW_c[14] , \BW_c[13] , \BW_c[12] , \BW_c[11] , \BW_c[10] , 
        \BW_c[9] , \BW_c[8] , \BW_c[7] , \BW_c[6] , \BW_c[5] , 
        \BW_c[4] , \BW_c[3] , \BW_c[2] , \BW_c[1] , \BW_c[0] }), 
        .dac1_db_c({\dac1_db_c[13] , \dac1_db_c[12] , \dac1_db_c[11] , 
        \dac1_db_c[10] , \dac1_db_c[9] , \dac1_db_c[8] , 
        \dac1_db_c[7] , \dac1_db_c[6] , \dac1_db_c[5] }), .temp1({
        \temp1[15] , \temp1[14] , \temp1[13] , \temp1[12] , 
        \temp1[11] , \temp1[10] , \temp1[9] , \temp1[8] , \temp1[7] , 
        \temp1[6] , \temp1[5] , \temp1[4] , \temp1[3] , \temp1[2] , 
        \temp1[1] , \temp1[0] }), .temp2({\temp2[15] , \temp2[14] , 
        \temp2[13] , \temp2[12] , \temp2[11] , \temp2[10] , \temp2[9] , 
        \temp2[8] , \temp2[7] , \temp2[6] , \temp2[5] , \temp2[4] , 
        \temp2[3] , \temp2[2] , \temp2[1] , \temp2[0] }), .temp3({
        \temp3[15] , \temp3[14] , \temp3[13] , \temp3[12] , 
        \temp3[11] , \temp3[10] , \temp3[9] , \temp3[8] , \temp3[7] , 
        \temp3[6] , \temp3[5] , \temp3[4] , \temp3[3] , \temp3[2] , 
        \temp3[1] , \temp3[0] }), .SENSE_DOUT_c({\SENSE_DOUT_c[1] }), 
        .temp_count({\temp_count[31] , \temp_count[30] , 
        \temp_count[29] , \temp_count[28] , \temp_count[27] , 
        \temp_count[26] , \temp_count[25] , \temp_count[24] , 
        \temp_count[23] , \temp_count[22] , \temp_count[21] , 
        \temp_count[20] , \temp_count[19] , \temp_count[18] , 
        \temp_count[17] , \temp_count[16] , \temp_count[15] , 
        \temp_count[14] , \temp_count[13] , \temp_count[12] , 
        \temp_count[11] , \temp_count[10] , \temp_count[9] , 
        \temp_count[8] , \temp_count[7] , \temp_count[6] , 
        \temp_count[5] , \temp_count[4] , \temp_count[3] , 
        \temp_count[2] , \temp_count[1] , \temp_count[0] }), .adc_d0_c({
        \adc_d0_c[13] , \adc_d0_c[12] , \adc_d0_c[11] , \adc_d0_c[10] , 
        \adc_d0_c[9] , \adc_d0_c[8] , \adc_d0_c[7] , \adc_d0_c[6] , 
        \adc_d0_c[5] , \adc_d0_c[4] , \adc_d0_c[3] , \adc_d0_c[2] , 
        \adc_d0_c[1] , \adc_d0_c[0] }), .freq_11(\freq[18] ), .freq_2(
        \freq[9] ), .freq_13(\freq[20] ), .freq_14(\freq[21] ), 
        .freq_15(\freq[22] ), .freq_0(\freq[7] ), .freq_1(\freq[8] ), 
        .freq_10(\freq[17] ), .freq_6(\freq[13] ), .GPIO20_c(GPIO20_c), 
        .temp_sck_c(temp_sck_c), .BW_clk_c(BW_clk_c), .BW_clk_c_i_0(
        BW_clk_c_i_0), .temp_so_c(temp_so_c), .GPIO4_c(GPIO4_c), 
        .temp_sck_c_i_0(temp_sck_c_i_0), .dac1_clk_c(dac1_clk_c), 
        .SENSE_CS_1_c(SENSE_CS_1_c), .GPIO16_c(GPIO16_c), .GPIO14_c(
        GPIO14_c), .GPIO7_c(GPIO7_c), .temp3_csn_c(temp3_csn_c), 
        .temp2_csn_c(temp2_csn_c), .temp1_csn_c(temp1_csn_c), 
        .GPIO11_c(GPIO11_c), .GPIO10_c(GPIO10_c), .dac2_clk_c(
        dac2_clk_c), .oclk_1_c(oclk_1_c), .osc_vcc_c(osc_vcc_c), 
        .adc_of_c(adc_of_c), .adc_oen_c(adc_oen_c), .adc_clk_c(
        adc_clk_c), .GPIO6_c(GPIO6_c), .ANTF_n2_c(ANTF_n2_c), 
        .ANTF_n1_c(ANTF_n1_c), .GPS1_LD_c(GPS1_LD_c), .GPS1_I1_c(
        GPS1_I1_c), .GPS1_I0_c(GPS1_I0_c), .GPIO9_c(GPIO9_c), 
        .GPS2_Q0_c(GPS2_Q0_c), .GPS2_LD_c(GPS2_LD_c), .GPS1_Q1_c(
        GPS1_Q1_c), .GPS1_Q0_c(GPS1_Q0_c), .GPS_I1_c(GPS_I1_c), 
        .GPS_I0_c(GPS_I0_c), .GPS2_Q1_c(GPS2_Q1_c), .GPIO3_c(GPIO3_c), 
        .GPIO5_c(GPIO5_c));
    TRIBUFF \fl_dq_obuft[7]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[7]));
    TRIBUFF \fl_dq_obuft[0]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[0]));
    OUTBUF \SENSE_DOUT_obuf[1]  (.D(\SENSE_DOUT_c[1] ), .PAD(
        SENSE_DOUT[1]));
    TRIBUFF sr_lbn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_lbn));
    TRIBUFF \fl_a_obuft[21]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[21]));
    INBUF ANTF_n1_ibuf (.PAD(ANTF_n1), .Y(ANTF_n1_c));
    INBUF \BW_ibuf[14]  (.PAD(BW[14]), .Y(\BW_c[14] ));
    OUTBUF adc_shdn_obuf (.D(VCC_net_1), .PAD(adc_shdn));
    TRIBUFF GPIO1_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(GPIO1));
    OUTBUF \dac1_db_obuf[9]  (.D(\dac1_db_c[9] ), .PAD(dac1_db[9]));
    OUTBUF \dac1_db_obuf[11]  (.D(\dac1_db_c[11] ), .PAD(dac1_db[11]));
    OUTBUF \dac1_db_obuf[6]  (.D(\dac1_db_c[6] ), .PAD(dac1_db[6]));
    TRIBUFF \fl_a_obuft[23]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[23]));
    OUTBUF CTR5_obuf (.D(GND_net_1), .PAD(CTR5));
    TRIBUFF \fl_dq_obuft[6]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[6]));
    TRIBUFF fl_cen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_cen));
    OUTBUF \dac1_db_obuf[10]  (.D(\dac1_db_c[10] ), .PAD(dac1_db[10]));
    INBUF \adc_d0_ibuf[13]  (.PAD(adc_d0[13]), .Y(\adc_d0_c[13] ));
    INBUF \BW_ibuf[2]  (.PAD(BW[2]), .Y(\BW_c[2] ));
    TRIBUFF REF_LE_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_LE));
    INBUF \BW_ibuf[11]  (.PAD(BW[11]), .Y(\BW_c[11] ));
    OUTBUF out1_obuf (.D(GND_net_1), .PAD(out1));
    OUTBUF CTR3_obuf (.D(GND_net_1), .PAD(CTR3));
    INBUF adc_oen_ibuf (.PAD(adc_oen), .Y(adc_oen_c));
    TRIBUFF REF_MXOUT_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        REF_MXOUT));
    INBUF \adc_d0_ibuf[9]  (.PAD(adc_d0[9]), .Y(\adc_d0_c[9] ));
    INBUF GPS1_I0_ibuf (.PAD(GPS1_I0), .Y(GPS1_I0_c));
    INBUF \adc_d0_ibuf[1]  (.PAD(adc_d0[1]), .Y(\adc_d0_c[1] ));
    TRIBUFF \fl_a_obuft[10]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[10]));
    OUTBUF CTR1_obuf (.D(GND_net_1), .PAD(CTR1));
    GND GND (.Y(GND_net_1));
    INBUF \SENSE_DIN_ibuf[0]  (.PAD(SENSE_DIN[0]), .Y(GPIO6_c));
    INBUF GPS2_Q0_ibuf (.PAD(GPS2_Q0), .Y(GPS2_Q0_c));
    OUTBUF \BW_out_obuf[11]  (.D(\BW_out_c[11] ), .PAD(BW_out[11]));
    OUTBUF \BW_out_obuf[6]  (.D(\BW_out_c[6] ), .PAD(BW_out[6]));
    OUTBUF \BW_out_obuf[1]  (.D(\BW_out_c[1] ), .PAD(BW_out[1]));
    OUTBUF GPIO12_obuf (.D(VCC_net_1), .PAD(GPIO12));
    OUTBUF GPIO15_obuf (.D(GND_net_1), .PAD(GPIO15));
    TRIBUFF \fl_a_obuft[17]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[17]));
    OUTBUF GPIO19_obuf (.D(GND_net_1), .PAD(GPIO19));
    TRIBUFF sr_cs2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_cs2));
    INBUF osc_vcc_ibuf (.PAD(osc_vcc), .Y(osc_vcc_c));
    syn_identify_core0_0 ident_coreinst (.temp1({\temp1[15] , 
        \temp1[14] , \temp1[13] , \temp1[12] , \temp1[11] , 
        \temp1[10] , \temp1[9] , \temp1[8] , \temp1[7] , \temp1[6] , 
        \temp1[5] , \temp1[4] , \temp1[3] , \temp1[2] , \temp1[1] , 
        \temp1[0] }), .temp2({\temp2[15] , \temp2[14] , \temp2[13] , 
        \temp2[12] , \temp2[11] , \temp2[10] , \temp2[9] , \temp2[8] , 
        \temp2[7] , \temp2[6] , \temp2[5] , \temp2[4] , \temp2[3] , 
        \temp2[2] , \temp2[1] , \temp2[0] }), .temp3({\temp3[15] , 
        \temp3[14] , \temp3[13] , \temp3[12] , \temp3[11] , 
        \temp3[10] , \temp3[9] , \temp3[8] , \temp3[7] , \temp3[6] , 
        \temp3[5] , \temp3[4] , \temp3[3] , \temp3[2] , \temp3[1] , 
        \temp3[0] }), .temp_count_data({\temp_count_data[4] , 
        \temp_count_data[3] , \temp_count_data[2] , 
        \temp_count_data[1] , \temp_count_data[0] }), .temp_count({
        \temp_count[31] , \temp_count[30] , \temp_count[29] , 
        \temp_count[28] , \temp_count[27] , \temp_count[26] , 
        \temp_count[25] , \temp_count[24] , \temp_count[23] , 
        \temp_count[22] , \temp_count[21] , \temp_count[20] , 
        \temp_count[19] , \temp_count[18] , \temp_count[17] , 
        \temp_count[16] , \temp_count[15] , \temp_count[14] , 
        \temp_count[13] , \temp_count[12] , \temp_count[11] , 
        \temp_count[10] , \temp_count[9] , \temp_count[8] , 
        \temp_count[7] , \temp_count[6] , \temp_count[5] , 
        \temp_count[4] , \temp_count[3] , \temp_count[2] , 
        \temp_count[1] , \temp_count[0] }), .freq_1(\freq[8] ), 
        .freq_2(\freq[9] ), .freq_0(\freq[7] ), .freq_6(\freq[13] ), 
        .freq_10(\freq[17] ), .freq_11(\freq[18] ), .freq_13(
        \freq[20] ), .freq_14(\freq[21] ), .freq_15(\freq[22] ), .atck(
        atck), .atdi(atdi), .atdo(atdo), .atms(atms), .atrstb(atrstb), 
        .BW_clk_c(BW_clk_c), .temp_sck_c(temp_sck_c), .temp1_csn_c(
        temp1_csn_c), .temp2_csn_c(temp2_csn_c), .temp3_csn_c(
        temp3_csn_c), .temp_so_c(temp_so_c));
    TRIBUFF dsa_le_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(dsa_le));
    INBUF \BW_ibuf[0]  (.PAD(BW[0]), .Y(\BW_c[0] ));
    TRIBUFF GPS1_SCLK_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_SCLK));
    TRIBUFF GPS1_PGM_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_PGM));
    TRIBUFF \fl_dq_obuft[3]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[3]));
    TRIBUFF \fl_a_obuft[12]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[12]));
    TRIBUFF GPS1_SHDN_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_SHDN));
    OUTBUF GPIO14_obuf (.D(GPIO14_c), .PAD(GPIO14));
    OUTBUF AMP_EN_obuf (.D(GND_net_1), .PAD(AMP_EN));
    INBUF \adc_d0_ibuf[3]  (.PAD(adc_d0[3]), .Y(\adc_d0_c[3] ));
    TRIBUFF \fl_a_obuft[15]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[15]));
    INBUF GPS1_Q1_ibuf (.PAD(GPS1_Q1), .Y(GPS1_Q1_c));
    OUTBUF \BW_out_obuf[10]  (.D(\BW_out_c[10] ), .PAD(BW_out[10]));
    TRIBUFF \SENSE_DOUT_obuft[0]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        SENSE_DOUT[0]));
    OUTBUF \BW_out_obuf[9]  (.D(\BW_out_c[9] ), .PAD(BW_out[9]));
    OUTBUF CTR4_obuf (.D(GND_net_1), .PAD(CTR4));
    VCC VCC (.Y(VCC_net_1));
    TRIBUFF fl_byten_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_byten));
    TRIBUFF \fl_a_obuft[0]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[0]));
    INBUF adc_clk_ibuf (.PAD(adc_clk), .Y(adc_clk_c));
    OUTBUF CTR2_obuf (.D(GND_net_1), .PAD(CTR2));
    TRIBUFF sr_ubn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_ubn));
    TRIBUFF dac1_sleep_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        dac1_sleep));
    TRIBUFF \fl_a_obuft[8]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[8]));
    TRIBUFF REF_CLK_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_CLK));
    TRIBUFF GPS1_IDLE_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_IDLE));
    TRIBUFF dsa_data_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        dsa_data));
    TRIBUFF en_modul_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        en_modul));
    INBUF \adc_d0_ibuf[11]  (.PAD(adc_d0[11]), .Y(\adc_d0_c[11] ));
    OUTBUF temp3_csn_obuf (.D(temp3_csn_c), .PAD(temp3_csn));
    TRIBUFF REF_DATA_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        REF_DATA));
    OUTBUF \dac1_db_obuf[8]  (.D(\dac1_db_c[8] ), .PAD(dac1_db[8]));
    TRIBUFF fl_oen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_oen));
    INBUF GPS1_LD_ibuf (.PAD(GPS1_LD), .Y(GPS1_LD_c));
    OUTBUF \dac1_db_obuf[5]  (.D(\dac1_db_c[5] ), .PAD(dac1_db[5]));
    INBUF \adc_d0_ibuf[10]  (.PAD(adc_d0[10]), .Y(\adc_d0_c[10] ));
    TRIBUFF \fl_a_obuft[20]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[20]));
    TRIBUFF CSN_n1_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(CSN_n1));
    INBUF GPS_I0_ibuf (.PAD(GPS_I0), .Y(GPS_I0_c));
    OUTBUF \BW_out_obuf[13]  (.D(\BW_out_c[13] ), .PAD(BW_out[13]));
    TRIBUFF \fl_a_obuft[4]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[4]));
    INBUF \adc_d0_ibuf[2]  (.PAD(adc_d0[2]), .Y(\adc_d0_c[2] ));
    OUTBUF CTR6_obuf (.D(GPIO8_c_i_0), .PAD(CTR6));
    INBUF GPS1_Q0_ibuf (.PAD(GPS1_Q0), .Y(GPS1_Q0_c));
    INBUF \BW_ibuf[6]  (.PAD(BW[6]), .Y(\BW_c[6] ));
    TRIBUFF \fl_dq_obuft[5]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[5]));
    CFG1 #( .INIT(2'h1) )  CTR7_obuf_RNO (.A(GPIO9_c), .Y(GPIO9_c_i_0));
    INBUF GPS2_LD_ibuf (.PAD(GPS2_LD), .Y(GPS2_LD_c));
    INBUF \BW_ibuf[10]  (.PAD(BW[10]), .Y(\BW_c[10] ));
    TRIBUFF fl_resetn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_resetn));
    OUTBUF \BW_out_obuf[12]  (.D(\BW_out_c[12] ), .PAD(BW_out[12]));
    OUTBUF GPIO6_obuf (.D(GPIO6_c), .PAD(GPIO6));
    TRIBUFF \fl_a_obuft[5]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[5]));
    TRIBUFF \fl_a_obuft[9]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[9]));
    CFG1 #( .INIT(2'h1) )  CTR6_obuf_RNO (.A(GPIO8_c), .Y(GPIO8_c_i_0));
    INBUF \BW_ibuf[8]  (.PAD(BW[8]), .Y(\BW_c[8] ));
    TRIBUFF fl_wen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_wen));
    TRIBUFF \fl_a_obuft[22]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[22]));
    TRIBUFF \fl_a_obuft[25]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[25]));
    OUTBUF BW_clk_obuf (.D(BW_clk_c), .PAD(BW_clk));
    TRIBUFF sr_oen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_oen));
    INBUF adc_of_ibuf (.PAD(adc_of), .Y(adc_of_c));
    INBUF GPIO9_ibuf (.PAD(GPIO9), .Y(GPIO9_c));
    INBUF GPIO8_ibuf (.PAD(GPIO8), .Y(GPIO8_c));
    TRIBUFF \fl_a_obuft[14]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[14]));
    TRIBUFF sr_wen_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_wen));
    INBUF \adc_d0_ibuf[4]  (.PAD(adc_d0[4]), .Y(\adc_d0_c[4] ));
    OUTBUF GPIO20_obuf (.D(GPIO20_c), .PAD(GPIO20));
    TRIBUFF BW_36_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(BW_36));
    TRIBUFF out2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(out2));
    OUTBUF \dac1_db_obuf[12]  (.D(\dac1_db_c[12] ), .PAD(dac1_db[12]));
    OUTBUF \BW_out_obuf[5]  (.D(\BW_out_c[5] ), .PAD(BW_out[5]));
    INBUF \BW_ibuf[12]  (.PAD(BW[12]), .Y(\BW_c[12] ));
    OUTBUF GPIO7_obuf (.D(GPIO7_c), .PAD(GPIO7));
    INBUF GPIO10_ibuf (.PAD(GPIO10), .Y(GPIO10_c));
    INBUF temp_so_ibuf (.PAD(temp_so), .Y(temp_so_c));
    TRIBUFF REF_CE_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_CE));
    INBUF \adc_d0_ibuf[0]  (.PAD(adc_d0[0]), .Y(\adc_d0_c[0] ));
    TRIBUFF \fl_a_obuft[18]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[18]));
    OUTBUF temp2_csn_obuf (.D(temp2_csn_c), .PAD(temp2_csn));
    OUTBUF CTR7_obuf (.D(GPIO9_c_i_0), .PAD(CTR7));
    TRIBUFF fl_wpn_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_wpn));
    INBUF \adc_d0_ibuf[5]  (.PAD(adc_d0[5]), .Y(\adc_d0_c[5] ));
    TRIBUFF dsa_clk_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(dsa_clk));
    TRIBUFF GPS1_SDATA_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        GPS1_SDATA));
    TRIBUFF \fl_dq_obuft[4]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[4]));
    OUTBUF \BW_out_obuf[14]  (.D(\BW_out_c[14] ), .PAD(BW_out[14]));
    OUTBUF \BW_out_obuf[0]  (.D(\BW_out_c[0] ), .PAD(BW_out[0]));
    TRIBUFF REF_LD_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(REF_LD));
    TRIBUFF clk_out_n2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        clk_out_n2));
    INBUF ANTF_n2_ibuf (.PAD(ANTF_n2), .Y(ANTF_n2_c));
    OUTBUF GPIO16_obuf (.D(GPIO16_c), .PAD(GPIO16));
    OUTBUF GPIO5_obuf (.D(GPIO5_c), .PAD(GPIO5));
    TRIBUFF \fl_a_obuft[11]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[11]));
    TRIBUFF \fl_a_obuft[19]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[19]));
    INBUF GPS_I1_ibuf (.PAD(GPS_I1), .Y(GPS_I1_c));
    TRIBUFF GPIO2_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(GPIO2));
    INBUF \SENSE_DIN_ibuf[1]  (.PAD(SENSE_DIN[1]), .Y(GPIO4_c));
    build_sb build_sb_0 (.temp_sck_c(temp_sck_c), .temp_sck_c_i_0(
        temp_sck_c_i_0), .BW_clk_c(BW_clk_c), .BW_clk_c_i_0(
        BW_clk_c_i_0));
    TRIBUFF \fl_a_obuft[6]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[6]));
    INBUF \BW_ibuf[7]  (.PAD(BW[7]), .Y(\BW_c[7] ));
    INBUF \adc_d0_ibuf[7]  (.PAD(adc_d0[7]), .Y(\adc_d0_c[7] ));
    TRIBUFF fl_ryby_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(fl_ryby));
    TRIBUFF \fl_a_obuft[13]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[13]));
    OUTBUF \dac1_db_obuf[7]  (.D(\dac1_db_c[7] ), .PAD(dac1_db[7]));
    OUTBUF GPIO4_obuf (.D(GPIO4_c), .PAD(GPIO4));
    OUTBUF temp1_csn_obuf (.D(temp1_csn_c), .PAD(temp1_csn));
    TRIBUFF \fl_a_obuft[1]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[1]));
    TRIBUFF \fl_a_obuft[3]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[3]));
    OUTBUF \dac1_db_obuf[13]  (.D(\dac1_db_c[13] ), .PAD(dac1_db[13]));
    TRIBUFF \fl_a_obuft[24]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[24]));
    INBUF \BW_ibuf[4]  (.PAD(BW[4]), .Y(\BW_c[4] ));
    INBUF \BW_ibuf[1]  (.PAD(BW[1]), .Y(\BW_c[1] ));
    OUTBUF temp_sck_obuf (.D(temp_sck_c), .PAD(temp_sck));
    TRIBUFF clk_out_n1_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(
        clk_out_n1));
    TRIBUFF \fl_a_obuft[16]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[16]));
    TRIBUFF \fl_dq_obuft[2]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_dq[2]));
    INBUF \BW_ibuf[13]  (.PAD(BW[13]), .Y(\BW_c[13] ));
    TRIBUFF \fl_a_obuft[7]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[7]));
    OUTBUF oclk_1_obuf (.D(oclk_1_c), .PAD(oclk_1));
    OUTBUF dac1_clk_obuf (.D(dac1_clk_c), .PAD(dac1_clk));
    OUTBUF \BW_out_obuf[2]  (.D(\BW_out_c[2] ), .PAD(BW_out[2]));
    TRIBUFF GPIO17_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(GPIO17));
    TRIBUFF sr_cs1n_obuft (.D(GND_net_1), .E(GND_net_1), .PAD(sr_cs1n));
    OUTBUF \BW_out_obuf[4]  (.D(\BW_out_c[4] ), .PAD(BW_out[4]));
    TRIBUFF \fl_a_obuft[2]  (.D(GND_net_1), .E(GND_net_1), .PAD(
        fl_a[2]));
    OUTBUF dac2_clk_obuf (.D(dac2_clk_c), .PAD(dac2_clk));
    OUTBUF SENSE_CS_1_obuf (.D(SENSE_CS_1_c), .PAD(SENSE_CS_1));
    INBUF GPIO11_ibuf (.PAD(GPIO11), .Y(GPIO11_c));
    INBUF \adc_d0_ibuf[12]  (.PAD(adc_d0[12]), .Y(\adc_d0_c[12] ));
    OUTBUF \BW_out_obuf[3]  (.D(\BW_out_c[3] ), .PAD(BW_out[3]));
    
endmodule
