// Target Device : IGLOO2 M2G010 484 FBGA
// Author : Malyshev
module led_igloo (
      input init_done,
      input fab_clk_100MHz,
      input fab_clk_8MHz,
      input fab_clk_5MHz,
      input fab_clk_1_17MHz,
      input temp_sck , // ???????????????? ?????????????? ????????????????????????????
      input temp_csn,  // ???????????????? ?????????????? ????????????????????????????
      input temp3_so,  // ???????????????? ?????????????? ????????????????????????????
      input temp2_so,  // ???????????????? ?????????????? ????????????????????????????
      input temp1_so,  // ???????????????? ?????????????? ????????????????????????????
      output reg out1,     // ???????????????? ??????????????????????
      output out2,     // ???????????????? ????????????????????????
      // ???????? ???????????????????? ????????????????
      input adc_clk,
      input [13:0] adc_d0,
      input adc_oen,
      input  adc_of,
      output reg adc_shdn = 1,

      input osc_vcc, // ???????????????????????? ???????????????????????????? ???????? GPS
      output reg [34:0] BW = 34'bz,   // ???????????????????????? ?????????????? ??????????
      output reg BW_36 = 0, // Reset neighbour FPGA
      // ???????? ?????????????????? ????????????????
      output dac1_clk,
      output dac2_clk,
      output reg [13:5] dac1_db,
      output dac1_sleep,
      // SRAM & FLASH
      output [25:0] fl_a,
      output fl_byten,
      output fl_cen,
      output [7:0] fl_dq,
      output fl_oen,
      output fl_resetn,
      output fl_ryby,
      output fl_wen,
      output fl_wpn,
      output sr_cs1n,
      output sr_cs2,
      output sr_lbn,
      output sr_oen,
      output sr_ubn,
      output sr_wen,
      // ???????????????????????????? GPS
      input ANTF_n1,
      output clk_out_n1,
      input  GPS1_I0,
      input GPS1_I1,
      input GPS1_LD,
      input GPS1_Q0,
      input GPS1_Q1,

      input ANTF_n2,
      output clk_out_n2,
      output CSN_n1,
      input GPS_I0,
      input GPS_I1,
      output GPS1_IDLE,
      input GPS2_LD,
      output GPS1_PGM,
      input GPS2_Q0,
      input GPS2_Q1,
      output GPS1_SCLK,
      output GPS1_SDATA,
      output GPS1_SHDN,
      // ???????????????????????????? ?????????????????????????????? ??????????????
      output REF_CE,
      output REF_CLK,
      output REF_DATA,
      output REF_LD,
      output REF_LE,
      output REF_MXOUT,
      // ???????? ???????? ???????? ????????????????????????????
      output reg SENSE_CS_1 = 1,
      input [1:0] SENSE_DIN,
      output reg [1:0] SENSE_DOUT,
      output oclk_1,
      // ???????????????????????????? ?????????????????????????????? ???????????????????? ????????????????
      output dsa_clk,
      output dsa_data,
      output dsa_le,
      // ???????????????????????? ????????????????????????
      output en_modul,
      output GPIO20,  //Den (RS485)
      output reg GPIO19 = 0,  // R (RS485)
      output GPIO17,  // SB3
      output reg GPIO16 = 1,  // LED3
      output reg GPIO15 = 0,  // D (RS485)
      output reg GPIO14 = 1,  // LED1
      output reg GPIO12,  // LED2
      input GPIO11,  // SB1
      input GPIO10,  // SB4
      input GPIO9,   // SB2
      input GPIO8,   // SB5
      output wire GPIO7,   // Ren (RS485)
      output wire GPIO6,
      output wire GPIO5,
      output wire GPIO4,
      output wire GPIO3,
      output GPIO2,   // RESETn
      output GPIO1,   // GOLDEN
      // ???????????????????????? ???????????????????????????????????? ???? 0.25 ????
      output reg CTR7 = 0,
      output reg CTR6 = 0,
      // *****
      output reg CTR5 = 0, // ???????????????????????? 0?? ???????? ??????????????????????????????
      output reg CTR4 = 0, // ???????????????????????? 0?? ???????? ??????????????????????
      output reg CTR3 = 0, // ???????????????????????? 5?? ???????? ??????????????????????????????
      output reg CTR2 = 0, // ???????????????????????? 5?? ???????? ??????????????????????
      output reg CTR1 = 0,  // ???????????????????????? 1?? ?????? ?????????????????????? ?????????????????????????????? ???????? ??????????????????????
      output reg AMP_EN = 0
  );

    reg [3:0] cnt_frame= 0;
    reg [9:0] cnt = 0;
    reg [31:0] freq;
    reg [31:0] cnt_freq = 0;
  
  assign GPIO5 = temp_sck^temp_csn^temp3_so^temp2_so^temp1_so^adc_clk^adc_oen^adc_of^osc_vcc^ANTF_n1^GPS1_I0^GPIO9^GPS1_I1^GPS1_LD^GPS1_Q0^GPS1_Q1^ANTF_n2^GPS_I0^GPS_I1^GPS2_LD^GPS2_Q0^GPS2_Q1^SENSE_DIN[0]^SENSE_DIN[1];
  assign GPIO6 = SENSE_DIN[0];
  assign GPIO4 = SENSE_DIN[1];
  assign GPIO7 = cnt[0]; 
  assign GPIO3 = adc_d0[13]^adc_d0[12]^adc_d0[11]^adc_d0[10]^adc_d0[9]^adc_d0[8]^adc_d0[7]^adc_d0[6]^adc_d0[5]^adc_d0[4]^adc_d0[3]^adc_d0[2]^adc_d0[1]^adc_d0[0];
  assign GPIO20 = SENSE_CS_1; 
  assign oclk_1 = fab_clk_8MHz*(~SENSE_CS_1); 


    reg [1:0] state = 2'b00;
    reg [7:0] data_2adc [8:0];
    reg [11:0] data_from_adc [8:0];
    
 
   always @ (posedge fab_clk_8MHz)
    begin
    data_2adc[0] = 8'b00_000_000; // none
    data_2adc[1] = 8'b11_000_111; // IN0
    data_2adc[2] = 8'b11_001_111; // IN1
    data_2adc[3] = 8'b11_010_111; // IN2
    data_2adc[4] = 8'b11_011_111; // IN3
    data_2adc[5] = 8'b11_100_111; // IN4
    data_2adc[6] = 8'b11_101_111; // IN5
    data_2adc[7] = 8'b11_110_111; // IN6
    data_2adc[8] = 8'b11_111_111; // IN7
    end
   
  always @ (negedge fab_clk_8MHz)
  begin
   case (state)
    2'b00 : begin
              if (!GPIO11)
               begin
                state <= 2'b01;
                cnt_frame <= 0;
               end
            end
    2'b01 : begin
             if (cnt_frame < 8)
                begin
                  cnt_frame <= cnt_frame + 1;
                  state <= 2'b10;
                  cnt <= 0; 
                end
             else
                state <= 2'b00;
            end
     2'b10 : begin
            if (cnt <=50)
            begin 
                cnt <= cnt + 1; 
             if (cnt <= 15 ) 
                    SENSE_CS_1 <= 0; 
             if (cnt >15 && cnt <= 50)
                    SENSE_CS_1 <= 1; 
             end 
             else 
                 begin
                    state <= 2'b01;
                    cnt <= 0;
                  end
              end 
     endcase
  end

    always @ (negedge fab_clk_8MHz) 
    begin 
         if (cnt > 0 && cnt <= 7)
            SENSE_DOUT[1] <= data_2adc[cnt_frame][7-cnt];
    end 

    always @ (posedge fab_clk_8MHz)
    begin 
        if (cnt >= 5 && cnt <= 16)
            data_from_adc [cnt_frame][16-cnt] <= SENSE_DIN[1];
    end 

    always @ (posedge fab_clk_8MHz)
    begin
       if ( $unsigned(data_from_adc[2][11:0]) < 12'd500 )
            freq <= 32'd400_000;
       if ( $unsigned(data_from_adc[2][11:0]) >= 12'd500 && $unsigned(data_from_adc[2][11:0]) < 12'd1500 )
            freq <= 32'd1_600_000;
       if ( $unsigned(data_from_adc[2][11:0]) >= 12'd1500 && $unsigned(data_from_adc[2][11:0]) < 12'd2500 )
            freq <= 32'd4_000_000;
        if ( $unsigned(data_from_adc[2][11:0]) >= 12'd2500 && $unsigned(data_from_adc[2][11:0]) < 12'd4095 )
            freq <= 32'd8_000_000;
    end

    always @ (posedge fab_clk_8MHz)
    begin
        if (cnt_freq < freq)
            cnt_freq <= cnt_freq + 1;
        else
            begin
            cnt_freq <= 0;
            GPIO16 <= ~GPIO16;
            end
        if (!init_done)
            GPIO12 <= 1;
    end
   
    
  endmodule
